`timescale 1ns/1ps

module xs_bugcase_tb (
    input  logic clock,
    input  logic reset,
    input  logic io_ctrl_ubtbEnable,
    input  logic io_ctrl_abtbEnable,
    input  logic io_ctrl_mbtbEnable,
    input  logic io_ctrl_tageEnable,
    input  logic io_ctrl_scEnable,
    input  logic io_ctrl_ittageEnable,
    input  logic [46:0] io_resetVector_addr,
    input  logic io_fromFtq_redirect_valid,
    input  logic [48:0] io_fromFtq_redirect_bits_cfiPc_addr,
    input  logic [48:0] io_fromFtq_redirect_bits_target_addr,
    input  logic io_fromFtq_redirect_bits_taken,
    input  logic [1:0] io_fromFtq_redirect_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_attribute_rasAction,
    input  logic io_fromFtq_redirect_bits_meta_phr_phrPtr_flag,
    input  logic [9:0] io_fromFtq_redirect_bits_meta_phr_phrPtr_value,
    input  logic [12:0] io_fromFtq_redirect_bits_meta_phr_phrLowBits,
    input  logic [15:0] io_fromFtq_redirect_bits_meta_commonHRMeta_ghr,
    input  logic [7:0] io_fromFtq_redirect_bits_meta_commonHRMeta_bw,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_0,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_1,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_2,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_3,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_4,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_5,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_6,
    input  logic io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_7,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_0_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_1_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_2_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_3_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_4_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_5_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_6_branchType,
    input  logic [1:0] io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_7_branchType,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_0,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_1,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_2,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_3,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_4,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_5,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_6,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_commonHRMeta_position_7,
    input  logic [3:0] io_fromFtq_redirect_bits_meta_ras_ssp,
    input  logic [2:0] io_fromFtq_redirect_bits_meta_ras_sctr,
    input  logic io_fromFtq_redirect_bits_meta_ras_tosw_flag,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_ras_tosw_value,
    input  logic io_fromFtq_redirect_bits_meta_ras_tosr_flag,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_ras_tosr_value,
    input  logic io_fromFtq_redirect_bits_meta_ras_nos_flag,
    input  logic [4:0] io_fromFtq_redirect_bits_meta_ras_nos_value,
    input  logic io_fromFtq_train_valid,
    input  logic [48:0] io_fromFtq_train_bits_startPc_addr,
    input  logic io_fromFtq_train_bits_branches_0_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_0_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_0_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_0_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_0_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_0_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_0_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_1_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_1_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_1_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_1_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_1_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_1_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_1_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_2_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_2_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_2_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_2_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_2_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_2_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_2_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_3_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_3_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_3_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_3_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_3_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_3_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_3_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_4_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_4_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_4_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_4_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_4_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_4_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_4_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_5_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_5_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_5_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_5_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_5_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_5_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_5_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_6_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_6_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_6_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_6_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_6_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_6_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_6_bits_mispredict,
    input  logic io_fromFtq_train_bits_branches_7_valid,
    input  logic [48:0] io_fromFtq_train_bits_branches_7_bits_target_addr,
    input  logic io_fromFtq_train_bits_branches_7_bits_taken,
    input  logic [4:0] io_fromFtq_train_bits_branches_7_bits_cfiPosition,
    input  logic [1:0] io_fromFtq_train_bits_branches_7_bits_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_branches_7_bits_attribute_rasAction,
    input  logic io_fromFtq_train_bits_branches_7_bits_mispredict,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_0_0_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_0_0_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_0_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_0_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_0_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_0_1_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_0_1_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_1_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_1_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_1_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_0_2_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_0_2_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_2_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_2_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_2_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_0_3_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_0_3_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_3_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_3_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_0_3_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_1_0_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_1_0_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_0_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_0_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_0_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_1_1_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_1_1_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_1_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_1_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_1_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_1_2_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_1_2_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_2_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_2_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_2_counter_value,
    input  logic io_fromFtq_train_bits_meta_mbtb_entries_1_3_rawHit,
    input  logic [4:0] io_fromFtq_train_bits_meta_mbtb_entries_1_3_position,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_3_attribute_branchType,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_3_attribute_rasAction,
    input  logic [1:0] io_fromFtq_train_bits_meta_mbtb_entries_1_3_counter_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_0_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_0_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_0_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_0_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_0_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_0_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_1_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_1_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_1_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_1_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_1_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_1_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_2_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_2_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_2_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_2_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_2_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_2_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_3_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_3_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_3_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_3_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_3_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_3_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_4_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_4_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_4_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_4_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_4_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_4_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_5_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_5_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_5_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_5_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_5_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_5_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_6_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_6_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_6_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_6_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_6_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_6_altOrBasePred,
    input  logic io_fromFtq_train_bits_meta_tage_entries_7_useProvider,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_7_providerTableIdx,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_7_providerWayIdx,
    input  logic [2:0] io_fromFtq_train_bits_meta_tage_entries_7_providerTakenCtr_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_tage_entries_7_providerUsefulCtr_value,
    input  logic io_fromFtq_train_bits_meta_tage_entries_7_altOrBasePred,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_0,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_1,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_2,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_3,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_4,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_5,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_6,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_0_7,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_0,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_1,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_2,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_3,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_4,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_5,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_6,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scPathResp_1_7,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_0,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_1,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_2,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_3,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_4,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_5,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_6,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_7,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_8,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_9,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_10,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_11,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_12,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_13,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_14,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_15,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_16,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_17,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_18,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_19,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_20,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_21,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_22,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_23,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_24,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_25,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_26,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_27,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_28,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_29,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_30,
    input  logic [5:0] io_fromFtq_train_bits_meta_sc_scBiasResp_31,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_0,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_1,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_2,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_3,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_4,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_5,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_6,
    input  logic [1:0] io_fromFtq_train_bits_meta_sc_scBiasLowerBits_7,
    input  logic io_fromFtq_train_bits_meta_sc_scCommonHR_valid,
    input  logic [15:0] io_fromFtq_train_bits_meta_sc_scCommonHR_ghr,
    input  logic [7:0] io_fromFtq_train_bits_meta_sc_scCommonHR_bw,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_0,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_1,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_2,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_3,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_4,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_5,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_6,
    input  logic io_fromFtq_train_bits_meta_sc_scPred_7,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_0,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_1,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_2,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_3,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_4,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_5,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_6,
    input  logic io_fromFtq_train_bits_meta_sc_tagePred_7,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_0,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_1,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_2,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_3,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_4,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_5,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_6,
    input  logic io_fromFtq_train_bits_meta_sc_tagePredValid_7,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_0,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_1,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_2,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_3,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_4,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_5,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_6,
    input  logic io_fromFtq_train_bits_meta_sc_useScPred_7,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_0,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_1,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_2,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_3,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_4,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_5,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_6,
    input  logic io_fromFtq_train_bits_meta_sc_sumAboveThres_7,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_0,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_1,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_2,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_3,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_4,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_5,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_6,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_7,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_0,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_1,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_2,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_3,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_4,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_5,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_6,
    input  logic io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_7,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predPathIdx_0,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predPathIdx_1,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predGlobalIdx_0,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predGlobalIdx_1,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predBWIdx_0,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predBWIdx_1,
    input  logic [6:0] io_fromFtq_train_bits_meta_sc_debug_predBiasIdx,
    input  logic io_fromFtq_train_bits_meta_ittage_provider_valid,
    input  logic [2:0] io_fromFtq_train_bits_meta_ittage_provider_bits,
    input  logic io_fromFtq_train_bits_meta_ittage_altProvider_valid,
    input  logic [2:0] io_fromFtq_train_bits_meta_ittage_altProvider_bits,
    input  logic io_fromFtq_train_bits_meta_ittage_altDiffers,
    input  logic io_fromFtq_train_bits_meta_ittage_providerUsefulCnt_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_ittage_providerCnt_value,
    input  logic [1:0] io_fromFtq_train_bits_meta_ittage_altProviderCnt_value,
    input  logic io_fromFtq_train_bits_meta_ittage_allocate_valid,
    input  logic [2:0] io_fromFtq_train_bits_meta_ittage_allocate_bits,
    input  logic [48:0] io_fromFtq_train_bits_meta_ittage_providerTarget_addr,
    input  logic [48:0] io_fromFtq_train_bits_meta_ittage_altProviderTarget_addr,
    input  logic [9:0] io_fromFtq_train_bits_meta_phr_phrPtr_value,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_phrLowBits,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_31_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_30_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_29_foldedHist,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_28_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_27_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_26_foldedHist,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_25_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_24_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_23_foldedHist,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_22_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_21_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_20_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_19_foldedHist,
    input  logic [7:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_18_foldedHist,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_17_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_16_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_15_foldedHist,
    input  logic [12:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_14_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_13_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_12_foldedHist,
    input  logic [11:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_11_foldedHist,
    input  logic [10:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_10_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_9_foldedHist,
    input  logic [7:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_8_foldedHist,
    input  logic [6:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_7_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_6_foldedHist,
    input  logic [7:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_5_foldedHist,
    input  logic [8:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_4_foldedHist,
    input  logic [7:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_3_foldedHist,
    input  logic [7:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_2_foldedHist,
    input  logic [6:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_1_foldedHist,
    input  logic [3:0] io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_0_foldedHist,
    input  logic io_fromFtq_commit_valid,
    input  logic [3:0] io_fromFtq_commit_bits_meta_ras_ssp,
    input  logic io_fromFtq_commit_bits_meta_ras_tosw_flag,
    input  logic [4:0] io_fromFtq_commit_bits_meta_ras_tosw_value,
    input  logic [1:0] io_fromFtq_commit_bits_attribute_rasAction,
    input  logic io_fromFtq_bpuPtr_flag,
    input  logic [5:0] io_fromFtq_bpuPtr_value,
    input  logic io_toFtq_prediction_ready,
    input  logic [7:0] boreChildrenBd_bore_array,
    input  logic boreChildrenBd_bore_all,
    input  logic boreChildrenBd_bore_req,
    input  logic boreChildrenBd_bore_writeen,
    input  logic [37:0] boreChildrenBd_bore_be,
    input  logic [9:0] boreChildrenBd_bore_addr,
    input  logic [111:0] boreChildrenBd_bore_indata,
    input  logic boreChildrenBd_bore_readen,
    input  logic [9:0] boreChildrenBd_bore_addr_rd,
    input  logic [7:0] boreChildrenBd_bore_1_array,
    input  logic boreChildrenBd_bore_1_all,
    input  logic boreChildrenBd_bore_1_req,
    input  logic boreChildrenBd_bore_1_writeen,
    input  logic [37:0] boreChildrenBd_bore_1_be,
    input  logic [7:0] boreChildrenBd_bore_1_addr,
    input  logic [37:0] boreChildrenBd_bore_1_indata,
    input  logic boreChildrenBd_bore_1_readen,
    input  logic [7:0] boreChildrenBd_bore_1_addr_rd,
    input  logic [7:0] boreChildrenBd_bore_2_array,
    input  logic boreChildrenBd_bore_2_all,
    input  logic boreChildrenBd_bore_2_req,
    input  logic boreChildrenBd_bore_2_writeen,
    input  logic [75:0] boreChildrenBd_bore_2_be,
    input  logic [7:0] boreChildrenBd_bore_2_addr,
    input  logic [75:0] boreChildrenBd_bore_2_indata,
    input  logic boreChildrenBd_bore_2_readen,
    input  logic [7:0] boreChildrenBd_bore_2_addr_rd,
    input  logic [7:0] boreChildrenBd_bore_3_array,
    input  logic boreChildrenBd_bore_3_all,
    input  logic boreChildrenBd_bore_3_req,
    input  logic boreChildrenBd_bore_3_writeen,
    input  logic [75:0] boreChildrenBd_bore_3_be,
    input  logic [7:0] boreChildrenBd_bore_3_addr,
    input  logic [75:0] boreChildrenBd_bore_3_indata,
    input  logic boreChildrenBd_bore_3_readen,
    input  logic [7:0] boreChildrenBd_bore_3_addr_rd,
    input  logic [7:0] boreChildrenBd_bore_4_array,
    input  logic boreChildrenBd_bore_4_all,
    input  logic boreChildrenBd_bore_4_req,
    input  logic boreChildrenBd_bore_4_writeen,
    input  logic [75:0] boreChildrenBd_bore_4_be,
    input  logic [7:0] boreChildrenBd_bore_4_addr,
    input  logic [75:0] boreChildrenBd_bore_4_indata,
    input  logic boreChildrenBd_bore_4_readen,
    input  logic [7:0] boreChildrenBd_bore_4_addr_rd,
    input  logic [7:0] boreChildrenBd_bore_5_addr,
    input  logic [7:0] boreChildrenBd_bore_5_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_5_wdata,
    input  logic [7:0] boreChildrenBd_bore_5_wmask,
    input  logic boreChildrenBd_bore_5_re,
    input  logic boreChildrenBd_bore_5_we,
    input  logic boreChildrenBd_bore_5_ack,
    input  logic boreChildrenBd_bore_5_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_5_array,
    input  logic [7:0] boreChildrenBd_bore_6_addr,
    input  logic [7:0] boreChildrenBd_bore_6_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_6_wdata,
    input  logic [7:0] boreChildrenBd_bore_6_wmask,
    input  logic boreChildrenBd_bore_6_re,
    input  logic boreChildrenBd_bore_6_we,
    input  logic boreChildrenBd_bore_6_ack,
    input  logic boreChildrenBd_bore_6_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_6_array,
    input  logic [7:0] boreChildrenBd_bore_7_addr,
    input  logic [7:0] boreChildrenBd_bore_7_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_7_wdata,
    input  logic [7:0] boreChildrenBd_bore_7_wmask,
    input  logic boreChildrenBd_bore_7_re,
    input  logic boreChildrenBd_bore_7_we,
    input  logic boreChildrenBd_bore_7_ack,
    input  logic boreChildrenBd_bore_7_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_7_array,
    input  logic [7:0] boreChildrenBd_bore_8_addr,
    input  logic [7:0] boreChildrenBd_bore_8_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_8_wdata,
    input  logic [7:0] boreChildrenBd_bore_8_wmask,
    input  logic boreChildrenBd_bore_8_re,
    input  logic boreChildrenBd_bore_8_we,
    input  logic boreChildrenBd_bore_8_ack,
    input  logic boreChildrenBd_bore_8_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_8_array,
    input  logic [7:0] boreChildrenBd_bore_9_addr,
    input  logic [7:0] boreChildrenBd_bore_9_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_9_wdata,
    input  logic [7:0] boreChildrenBd_bore_9_wmask,
    input  logic boreChildrenBd_bore_9_re,
    input  logic boreChildrenBd_bore_9_we,
    input  logic boreChildrenBd_bore_9_ack,
    input  logic boreChildrenBd_bore_9_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_9_array,
    input  logic [7:0] boreChildrenBd_bore_10_addr,
    input  logic [7:0] boreChildrenBd_bore_10_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_10_wdata,
    input  logic [7:0] boreChildrenBd_bore_10_wmask,
    input  logic boreChildrenBd_bore_10_re,
    input  logic boreChildrenBd_bore_10_we,
    input  logic boreChildrenBd_bore_10_ack,
    input  logic boreChildrenBd_bore_10_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_10_array,
    input  logic [7:0] boreChildrenBd_bore_11_addr,
    input  logic [7:0] boreChildrenBd_bore_11_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_11_wdata,
    input  logic [7:0] boreChildrenBd_bore_11_wmask,
    input  logic boreChildrenBd_bore_11_re,
    input  logic boreChildrenBd_bore_11_we,
    input  logic boreChildrenBd_bore_11_ack,
    input  logic boreChildrenBd_bore_11_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_11_array,
    input  logic [7:0] boreChildrenBd_bore_12_addr,
    input  logic [7:0] boreChildrenBd_bore_12_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_12_wdata,
    input  logic [7:0] boreChildrenBd_bore_12_wmask,
    input  logic boreChildrenBd_bore_12_re,
    input  logic boreChildrenBd_bore_12_we,
    input  logic boreChildrenBd_bore_12_ack,
    input  logic boreChildrenBd_bore_12_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_12_array,
    input  logic [7:0] boreChildrenBd_bore_13_addr,
    input  logic [7:0] boreChildrenBd_bore_13_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_13_wdata,
    input  logic [7:0] boreChildrenBd_bore_13_wmask,
    input  logic boreChildrenBd_bore_13_re,
    input  logic boreChildrenBd_bore_13_we,
    input  logic boreChildrenBd_bore_13_ack,
    input  logic boreChildrenBd_bore_13_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_13_array,
    input  logic [7:0] boreChildrenBd_bore_14_addr,
    input  logic [7:0] boreChildrenBd_bore_14_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_14_wdata,
    input  logic [7:0] boreChildrenBd_bore_14_wmask,
    input  logic boreChildrenBd_bore_14_re,
    input  logic boreChildrenBd_bore_14_we,
    input  logic boreChildrenBd_bore_14_ack,
    input  logic boreChildrenBd_bore_14_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_14_array,
    input  logic [7:0] boreChildrenBd_bore_15_addr,
    input  logic [7:0] boreChildrenBd_bore_15_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_15_wdata,
    input  logic [7:0] boreChildrenBd_bore_15_wmask,
    input  logic boreChildrenBd_bore_15_re,
    input  logic boreChildrenBd_bore_15_we,
    input  logic boreChildrenBd_bore_15_ack,
    input  logic boreChildrenBd_bore_15_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_15_array,
    input  logic [7:0] boreChildrenBd_bore_16_addr,
    input  logic [7:0] boreChildrenBd_bore_16_addr_rd,
    input  logic [47:0] boreChildrenBd_bore_16_wdata,
    input  logic [7:0] boreChildrenBd_bore_16_wmask,
    input  logic boreChildrenBd_bore_16_re,
    input  logic boreChildrenBd_bore_16_we,
    input  logic boreChildrenBd_bore_16_ack,
    input  logic boreChildrenBd_bore_16_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_16_array,
    input  logic [7:0] boreChildrenBd_bore_17_addr,
    input  logic [7:0] boreChildrenBd_bore_17_addr_rd,
    input  logic [191:0] boreChildrenBd_bore_17_wdata,
    input  logic [31:0] boreChildrenBd_bore_17_wmask,
    input  logic boreChildrenBd_bore_17_re,
    input  logic boreChildrenBd_bore_17_we,
    input  logic boreChildrenBd_bore_17_ack,
    input  logic boreChildrenBd_bore_17_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_17_array,
    input  logic [7:0] boreChildrenBd_bore_18_addr,
    input  logic [7:0] boreChildrenBd_bore_18_addr_rd,
    input  logic [191:0] boreChildrenBd_bore_18_wdata,
    input  logic [31:0] boreChildrenBd_bore_18_wmask,
    input  logic boreChildrenBd_bore_18_re,
    input  logic boreChildrenBd_bore_18_we,
    input  logic boreChildrenBd_bore_18_ack,
    input  logic boreChildrenBd_bore_18_selectedOH,
    input  logic [7:0] boreChildrenBd_bore_18_array,
    input  logic sigFromSrams_bore_ram_hold,
    input  logic sigFromSrams_bore_ram_bypass,
    input  logic sigFromSrams_bore_ram_bp_clken,
    input  logic sigFromSrams_bore_ram_aux_clk,
    input  logic sigFromSrams_bore_ram_aux_ckbp,
    input  logic sigFromSrams_bore_ram_mcp_hold,
    input  logic sigFromSrams_bore_cgen,
    input  logic sigFromSrams_bore_1_ram_hold,
    input  logic sigFromSrams_bore_1_ram_bypass,
    input  logic sigFromSrams_bore_1_ram_bp_clken,
    input  logic sigFromSrams_bore_1_ram_aux_clk,
    input  logic sigFromSrams_bore_1_ram_aux_ckbp,
    input  logic sigFromSrams_bore_1_ram_mcp_hold,
    input  logic sigFromSrams_bore_1_cgen,
    input  logic sigFromSrams_bore_2_ram_hold,
    input  logic sigFromSrams_bore_2_ram_bypass,
    input  logic sigFromSrams_bore_2_ram_bp_clken,
    input  logic sigFromSrams_bore_2_ram_aux_clk,
    input  logic sigFromSrams_bore_2_ram_aux_ckbp,
    input  logic sigFromSrams_bore_2_ram_mcp_hold,
    input  logic sigFromSrams_bore_2_cgen,
    input  logic sigFromSrams_bore_3_ram_hold,
    input  logic sigFromSrams_bore_3_ram_bypass,
    input  logic sigFromSrams_bore_3_ram_bp_clken,
    input  logic sigFromSrams_bore_3_ram_aux_clk,
    input  logic sigFromSrams_bore_3_ram_aux_ckbp,
    input  logic sigFromSrams_bore_3_ram_mcp_hold,
    input  logic sigFromSrams_bore_3_cgen,
    input  logic sigFromSrams_bore_4_ram_hold,
    input  logic sigFromSrams_bore_4_ram_bypass,
    input  logic sigFromSrams_bore_4_ram_bp_clken,
    input  logic sigFromSrams_bore_4_ram_aux_clk,
    input  logic sigFromSrams_bore_4_ram_aux_ckbp,
    input  logic sigFromSrams_bore_4_ram_mcp_hold,
    input  logic sigFromSrams_bore_4_cgen,
    input  logic sigFromSrams_bore_5_ram_hold,
    input  logic sigFromSrams_bore_5_ram_bypass,
    input  logic sigFromSrams_bore_5_ram_bp_clken,
    input  logic sigFromSrams_bore_5_ram_aux_clk,
    input  logic sigFromSrams_bore_5_ram_aux_ckbp,
    input  logic sigFromSrams_bore_5_ram_mcp_hold,
    input  logic sigFromSrams_bore_5_cgen,
    input  logic sigFromSrams_bore_6_ram_hold,
    input  logic sigFromSrams_bore_6_ram_bypass,
    input  logic sigFromSrams_bore_6_ram_bp_clken,
    input  logic sigFromSrams_bore_6_ram_aux_clk,
    input  logic sigFromSrams_bore_6_ram_aux_ckbp,
    input  logic sigFromSrams_bore_6_ram_mcp_hold,
    input  logic sigFromSrams_bore_6_cgen,
    input  logic sigFromSrams_bore_7_ram_hold,
    input  logic sigFromSrams_bore_7_ram_bypass,
    input  logic sigFromSrams_bore_7_ram_bp_clken,
    input  logic sigFromSrams_bore_7_ram_aux_clk,
    input  logic sigFromSrams_bore_7_ram_aux_ckbp,
    input  logic sigFromSrams_bore_7_ram_mcp_hold,
    input  logic sigFromSrams_bore_7_cgen,
    input  logic sigFromSrams_bore_8_ram_hold,
    input  logic sigFromSrams_bore_8_ram_bypass,
    input  logic sigFromSrams_bore_8_ram_bp_clken,
    input  logic sigFromSrams_bore_8_ram_aux_clk,
    input  logic sigFromSrams_bore_8_ram_aux_ckbp,
    input  logic sigFromSrams_bore_8_ram_mcp_hold,
    input  logic sigFromSrams_bore_8_cgen,
    input  logic sigFromSrams_bore_9_ram_hold,
    input  logic sigFromSrams_bore_9_ram_bypass,
    input  logic sigFromSrams_bore_9_ram_bp_clken,
    input  logic sigFromSrams_bore_9_ram_aux_clk,
    input  logic sigFromSrams_bore_9_ram_aux_ckbp,
    input  logic sigFromSrams_bore_9_ram_mcp_hold,
    input  logic sigFromSrams_bore_9_cgen,
    input  logic sigFromSrams_bore_10_ram_hold,
    input  logic sigFromSrams_bore_10_ram_bypass,
    input  logic sigFromSrams_bore_10_ram_bp_clken,
    input  logic sigFromSrams_bore_10_ram_aux_clk,
    input  logic sigFromSrams_bore_10_ram_aux_ckbp,
    input  logic sigFromSrams_bore_10_ram_mcp_hold,
    input  logic sigFromSrams_bore_10_cgen,
    input  logic sigFromSrams_bore_11_ram_hold,
    input  logic sigFromSrams_bore_11_ram_bypass,
    input  logic sigFromSrams_bore_11_ram_bp_clken,
    input  logic sigFromSrams_bore_11_ram_aux_clk,
    input  logic sigFromSrams_bore_11_ram_aux_ckbp,
    input  logic sigFromSrams_bore_11_ram_mcp_hold,
    input  logic sigFromSrams_bore_11_cgen,
    input  logic sigFromSrams_bore_12_ram_hold,
    input  logic sigFromSrams_bore_12_ram_bypass,
    input  logic sigFromSrams_bore_12_ram_bp_clken,
    input  logic sigFromSrams_bore_12_ram_aux_clk,
    input  logic sigFromSrams_bore_12_ram_aux_ckbp,
    input  logic sigFromSrams_bore_12_ram_mcp_hold,
    input  logic sigFromSrams_bore_12_cgen,
    input  logic sigFromSrams_bore_13_ram_hold,
    input  logic sigFromSrams_bore_13_ram_bypass,
    input  logic sigFromSrams_bore_13_ram_bp_clken,
    input  logic sigFromSrams_bore_13_ram_aux_clk,
    input  logic sigFromSrams_bore_13_ram_aux_ckbp,
    input  logic sigFromSrams_bore_13_ram_mcp_hold,
    input  logic sigFromSrams_bore_13_cgen,
    input  logic sigFromSrams_bore_14_ram_hold,
    input  logic sigFromSrams_bore_14_ram_bypass,
    input  logic sigFromSrams_bore_14_ram_bp_clken,
    input  logic sigFromSrams_bore_14_ram_aux_clk,
    input  logic sigFromSrams_bore_14_ram_aux_ckbp,
    input  logic sigFromSrams_bore_14_ram_mcp_hold,
    input  logic sigFromSrams_bore_14_cgen,
    input  logic sigFromSrams_bore_15_ram_hold,
    input  logic sigFromSrams_bore_15_ram_bypass,
    input  logic sigFromSrams_bore_15_ram_bp_clken,
    input  logic sigFromSrams_bore_15_ram_aux_clk,
    input  logic sigFromSrams_bore_15_ram_aux_ckbp,
    input  logic sigFromSrams_bore_15_ram_mcp_hold,
    input  logic sigFromSrams_bore_15_cgen,
    input  logic sigFromSrams_bore_16_ram_hold,
    input  logic sigFromSrams_bore_16_ram_bypass,
    input  logic sigFromSrams_bore_16_ram_bp_clken,
    input  logic sigFromSrams_bore_16_ram_aux_clk,
    input  logic sigFromSrams_bore_16_ram_aux_ckbp,
    input  logic sigFromSrams_bore_16_ram_mcp_hold,
    input  logic sigFromSrams_bore_16_cgen,
    input  logic sigFromSrams_bore_17_ram_hold,
    input  logic sigFromSrams_bore_17_ram_bypass,
    input  logic sigFromSrams_bore_17_ram_bp_clken,
    input  logic sigFromSrams_bore_17_ram_aux_clk,
    input  logic sigFromSrams_bore_17_ram_aux_ckbp,
    input  logic sigFromSrams_bore_17_ram_mcp_hold,
    input  logic sigFromSrams_bore_17_cgen,
    input  logic sigFromSrams_bore_18_ram_hold,
    input  logic sigFromSrams_bore_18_ram_bypass,
    input  logic sigFromSrams_bore_18_ram_bp_clken,
    input  logic sigFromSrams_bore_18_ram_aux_clk,
    input  logic sigFromSrams_bore_18_ram_aux_ckbp,
    input  logic sigFromSrams_bore_18_ram_mcp_hold,
    input  logic sigFromSrams_bore_18_cgen,
    input  logic sigFromSrams_bore_19_ram_hold,
    input  logic sigFromSrams_bore_19_ram_bypass,
    input  logic sigFromSrams_bore_19_ram_bp_clken,
    input  logic sigFromSrams_bore_19_ram_aux_clk,
    input  logic sigFromSrams_bore_19_ram_aux_ckbp,
    input  logic sigFromSrams_bore_19_ram_mcp_hold,
    input  logic sigFromSrams_bore_19_cgen,
    input  logic sigFromSrams_bore_20_ram_hold,
    input  logic sigFromSrams_bore_20_ram_bypass,
    input  logic sigFromSrams_bore_20_ram_bp_clken,
    input  logic sigFromSrams_bore_20_ram_aux_clk,
    input  logic sigFromSrams_bore_20_ram_aux_ckbp,
    input  logic sigFromSrams_bore_20_ram_mcp_hold,
    input  logic sigFromSrams_bore_20_cgen,
    input  logic sigFromSrams_bore_21_ram_hold,
    input  logic sigFromSrams_bore_21_ram_bypass,
    input  logic sigFromSrams_bore_21_ram_bp_clken,
    input  logic sigFromSrams_bore_21_ram_aux_clk,
    input  logic sigFromSrams_bore_21_ram_aux_ckbp,
    input  logic sigFromSrams_bore_21_ram_mcp_hold,
    input  logic sigFromSrams_bore_21_cgen,
    input  logic sigFromSrams_bore_22_ram_hold,
    input  logic sigFromSrams_bore_22_ram_bypass,
    input  logic sigFromSrams_bore_22_ram_bp_clken,
    input  logic sigFromSrams_bore_22_ram_aux_clk,
    input  logic sigFromSrams_bore_22_ram_aux_ckbp,
    input  logic sigFromSrams_bore_22_ram_mcp_hold,
    input  logic sigFromSrams_bore_22_cgen,
    input  logic sigFromSrams_bore_23_ram_hold,
    input  logic sigFromSrams_bore_23_ram_bypass,
    input  logic sigFromSrams_bore_23_ram_bp_clken,
    input  logic sigFromSrams_bore_23_ram_aux_clk,
    input  logic sigFromSrams_bore_23_ram_aux_ckbp,
    input  logic sigFromSrams_bore_23_ram_mcp_hold,
    input  logic sigFromSrams_bore_23_cgen,
    input  logic sigFromSrams_bore_24_ram_hold,
    input  logic sigFromSrams_bore_24_ram_bypass,
    input  logic sigFromSrams_bore_24_ram_bp_clken,
    input  logic sigFromSrams_bore_24_ram_aux_clk,
    input  logic sigFromSrams_bore_24_ram_aux_ckbp,
    input  logic sigFromSrams_bore_24_ram_mcp_hold,
    input  logic sigFromSrams_bore_24_cgen,
    input  logic sigFromSrams_bore_25_ram_hold,
    input  logic sigFromSrams_bore_25_ram_bypass,
    input  logic sigFromSrams_bore_25_ram_bp_clken,
    input  logic sigFromSrams_bore_25_ram_aux_clk,
    input  logic sigFromSrams_bore_25_ram_aux_ckbp,
    input  logic sigFromSrams_bore_25_ram_mcp_hold,
    input  logic sigFromSrams_bore_25_cgen,
    input  logic sigFromSrams_bore_26_ram_hold,
    input  logic sigFromSrams_bore_26_ram_bypass,
    input  logic sigFromSrams_bore_26_ram_bp_clken,
    input  logic sigFromSrams_bore_26_ram_aux_clk,
    input  logic sigFromSrams_bore_26_ram_aux_ckbp,
    input  logic sigFromSrams_bore_26_ram_mcp_hold,
    input  logic sigFromSrams_bore_26_cgen,
    input  logic sigFromSrams_bore_27_ram_hold,
    input  logic sigFromSrams_bore_27_ram_bypass,
    input  logic sigFromSrams_bore_27_ram_bp_clken,
    input  logic sigFromSrams_bore_27_ram_aux_clk,
    input  logic sigFromSrams_bore_27_ram_aux_ckbp,
    input  logic sigFromSrams_bore_27_ram_mcp_hold,
    input  logic sigFromSrams_bore_27_cgen,
    input  logic sigFromSrams_bore_28_ram_hold,
    input  logic sigFromSrams_bore_28_ram_bypass,
    input  logic sigFromSrams_bore_28_ram_bp_clken,
    input  logic sigFromSrams_bore_28_ram_aux_clk,
    input  logic sigFromSrams_bore_28_ram_aux_ckbp,
    input  logic sigFromSrams_bore_28_ram_mcp_hold,
    input  logic sigFromSrams_bore_28_cgen,
    input  logic sigFromSrams_bore_29_ram_hold,
    input  logic sigFromSrams_bore_29_ram_bypass,
    input  logic sigFromSrams_bore_29_ram_bp_clken,
    input  logic sigFromSrams_bore_29_ram_aux_clk,
    input  logic sigFromSrams_bore_29_ram_aux_ckbp,
    input  logic sigFromSrams_bore_29_ram_mcp_hold,
    input  logic sigFromSrams_bore_29_cgen,
    input  logic sigFromSrams_bore_30_ram_hold,
    input  logic sigFromSrams_bore_30_ram_bypass,
    input  logic sigFromSrams_bore_30_ram_bp_clken,
    input  logic sigFromSrams_bore_30_ram_aux_clk,
    input  logic sigFromSrams_bore_30_ram_aux_ckbp,
    input  logic sigFromSrams_bore_30_ram_mcp_hold,
    input  logic sigFromSrams_bore_30_cgen,
    input  logic sigFromSrams_bore_31_ram_hold,
    input  logic sigFromSrams_bore_31_ram_bypass,
    input  logic sigFromSrams_bore_31_ram_bp_clken,
    input  logic sigFromSrams_bore_31_ram_aux_clk,
    input  logic sigFromSrams_bore_31_ram_aux_ckbp,
    input  logic sigFromSrams_bore_31_ram_mcp_hold,
    input  logic sigFromSrams_bore_31_cgen,
    input  logic sigFromSrams_bore_32_ram_hold,
    input  logic sigFromSrams_bore_32_ram_bypass,
    input  logic sigFromSrams_bore_32_ram_bp_clken,
    input  logic sigFromSrams_bore_32_ram_aux_clk,
    input  logic sigFromSrams_bore_32_ram_aux_ckbp,
    input  logic sigFromSrams_bore_32_ram_mcp_hold,
    input  logic sigFromSrams_bore_32_cgen,
    input  logic sigFromSrams_bore_33_ram_hold,
    input  logic sigFromSrams_bore_33_ram_bypass,
    input  logic sigFromSrams_bore_33_ram_bp_clken,
    input  logic sigFromSrams_bore_33_ram_aux_clk,
    input  logic sigFromSrams_bore_33_ram_aux_ckbp,
    input  logic sigFromSrams_bore_33_ram_mcp_hold,
    input  logic sigFromSrams_bore_33_cgen,
    input  logic sigFromSrams_bore_34_ram_hold,
    input  logic sigFromSrams_bore_34_ram_bypass,
    input  logic sigFromSrams_bore_34_ram_bp_clken,
    input  logic sigFromSrams_bore_34_ram_aux_clk,
    input  logic sigFromSrams_bore_34_ram_aux_ckbp,
    input  logic sigFromSrams_bore_34_ram_mcp_hold,
    input  logic sigFromSrams_bore_34_cgen,
    input  logic sigFromSrams_bore_35_ram_hold,
    input  logic sigFromSrams_bore_35_ram_bypass,
    input  logic sigFromSrams_bore_35_ram_bp_clken,
    input  logic sigFromSrams_bore_35_ram_aux_clk,
    input  logic sigFromSrams_bore_35_ram_aux_ckbp,
    input  logic sigFromSrams_bore_35_ram_mcp_hold,
    input  logic sigFromSrams_bore_35_cgen,
    input  logic sigFromSrams_bore_36_ram_hold,
    input  logic sigFromSrams_bore_36_ram_bypass,
    input  logic sigFromSrams_bore_36_ram_bp_clken,
    input  logic sigFromSrams_bore_36_ram_aux_clk,
    input  logic sigFromSrams_bore_36_ram_aux_ckbp,
    input  logic sigFromSrams_bore_36_ram_mcp_hold,
    input  logic sigFromSrams_bore_36_cgen,
    input  logic sigFromSrams_bore_37_ram_hold,
    input  logic sigFromSrams_bore_37_ram_bypass,
    input  logic sigFromSrams_bore_37_ram_bp_clken,
    input  logic sigFromSrams_bore_37_ram_aux_clk,
    input  logic sigFromSrams_bore_37_ram_aux_ckbp,
    input  logic sigFromSrams_bore_37_ram_mcp_hold,
    input  logic sigFromSrams_bore_37_cgen,
    input  logic sigFromSrams_bore_38_ram_hold,
    input  logic sigFromSrams_bore_38_ram_bypass,
    input  logic sigFromSrams_bore_38_ram_bp_clken,
    input  logic sigFromSrams_bore_38_ram_aux_clk,
    input  logic sigFromSrams_bore_38_ram_aux_ckbp,
    input  logic sigFromSrams_bore_38_ram_mcp_hold,
    input  logic sigFromSrams_bore_38_cgen,
    input  logic sigFromSrams_bore_39_ram_hold,
    input  logic sigFromSrams_bore_39_ram_bypass,
    input  logic sigFromSrams_bore_39_ram_bp_clken,
    input  logic sigFromSrams_bore_39_ram_aux_clk,
    input  logic sigFromSrams_bore_39_ram_aux_ckbp,
    input  logic sigFromSrams_bore_39_ram_mcp_hold,
    input  logic sigFromSrams_bore_39_cgen,
    input  logic sigFromSrams_bore_40_ram_hold,
    input  logic sigFromSrams_bore_40_ram_bypass,
    input  logic sigFromSrams_bore_40_ram_bp_clken,
    input  logic sigFromSrams_bore_40_ram_aux_clk,
    input  logic sigFromSrams_bore_40_ram_aux_ckbp,
    input  logic sigFromSrams_bore_40_ram_mcp_hold,
    input  logic sigFromSrams_bore_40_cgen,
    input  logic sigFromSrams_bore_41_ram_hold,
    input  logic sigFromSrams_bore_41_ram_bypass,
    input  logic sigFromSrams_bore_41_ram_bp_clken,
    input  logic sigFromSrams_bore_41_ram_aux_clk,
    input  logic sigFromSrams_bore_41_ram_aux_ckbp,
    input  logic sigFromSrams_bore_41_ram_mcp_hold,
    input  logic sigFromSrams_bore_41_cgen,
    input  logic sigFromSrams_bore_42_ram_hold,
    input  logic sigFromSrams_bore_42_ram_bypass,
    input  logic sigFromSrams_bore_42_ram_bp_clken,
    input  logic sigFromSrams_bore_42_ram_aux_clk,
    input  logic sigFromSrams_bore_42_ram_aux_ckbp,
    input  logic sigFromSrams_bore_42_ram_mcp_hold,
    input  logic sigFromSrams_bore_42_cgen,
    input  logic sigFromSrams_bore_43_ram_hold,
    input  logic sigFromSrams_bore_43_ram_bypass,
    input  logic sigFromSrams_bore_43_ram_bp_clken,
    input  logic sigFromSrams_bore_43_ram_aux_clk,
    input  logic sigFromSrams_bore_43_ram_aux_ckbp,
    input  logic sigFromSrams_bore_43_ram_mcp_hold,
    input  logic sigFromSrams_bore_43_cgen,
    input  logic sigFromSrams_bore_44_ram_hold,
    input  logic sigFromSrams_bore_44_ram_bypass,
    input  logic sigFromSrams_bore_44_ram_bp_clken,
    input  logic sigFromSrams_bore_44_ram_aux_clk,
    input  logic sigFromSrams_bore_44_ram_aux_ckbp,
    input  logic sigFromSrams_bore_44_ram_mcp_hold,
    input  logic sigFromSrams_bore_44_cgen,
    input  logic sigFromSrams_bore_45_ram_hold,
    input  logic sigFromSrams_bore_45_ram_bypass,
    input  logic sigFromSrams_bore_45_ram_bp_clken,
    input  logic sigFromSrams_bore_45_ram_aux_clk,
    input  logic sigFromSrams_bore_45_ram_aux_ckbp,
    input  logic sigFromSrams_bore_45_ram_mcp_hold,
    input  logic sigFromSrams_bore_45_cgen,
    input  logic sigFromSrams_bore_46_ram_hold,
    input  logic sigFromSrams_bore_46_ram_bypass,
    input  logic sigFromSrams_bore_46_ram_bp_clken,
    input  logic sigFromSrams_bore_46_ram_aux_clk,
    input  logic sigFromSrams_bore_46_ram_aux_ckbp,
    input  logic sigFromSrams_bore_46_ram_mcp_hold,
    input  logic sigFromSrams_bore_46_cgen,
    input  logic sigFromSrams_bore_47_ram_hold,
    input  logic sigFromSrams_bore_47_ram_bypass,
    input  logic sigFromSrams_bore_47_ram_bp_clken,
    input  logic sigFromSrams_bore_47_ram_aux_clk,
    input  logic sigFromSrams_bore_47_ram_aux_ckbp,
    input  logic sigFromSrams_bore_47_ram_mcp_hold,
    input  logic sigFromSrams_bore_47_cgen,
    input  logic sigFromSrams_bore_48_ram_hold,
    input  logic sigFromSrams_bore_48_ram_bypass,
    input  logic sigFromSrams_bore_48_ram_bp_clken,
    input  logic sigFromSrams_bore_48_ram_aux_clk,
    input  logic sigFromSrams_bore_48_ram_aux_ckbp,
    input  logic sigFromSrams_bore_48_ram_mcp_hold,
    input  logic sigFromSrams_bore_48_cgen,
    input  logic sigFromSrams_bore_49_ram_hold,
    input  logic sigFromSrams_bore_49_ram_bypass,
    input  logic sigFromSrams_bore_49_ram_bp_clken,
    input  logic sigFromSrams_bore_49_ram_aux_clk,
    input  logic sigFromSrams_bore_49_ram_aux_ckbp,
    input  logic sigFromSrams_bore_49_ram_mcp_hold,
    input  logic sigFromSrams_bore_49_cgen,
    input  logic sigFromSrams_bore_50_ram_hold,
    input  logic sigFromSrams_bore_50_ram_bypass,
    input  logic sigFromSrams_bore_50_ram_bp_clken,
    input  logic sigFromSrams_bore_50_ram_aux_clk,
    input  logic sigFromSrams_bore_50_ram_aux_ckbp,
    input  logic sigFromSrams_bore_50_ram_mcp_hold,
    input  logic sigFromSrams_bore_50_cgen,
    input  logic sigFromSrams_bore_51_ram_hold,
    input  logic sigFromSrams_bore_51_ram_bypass,
    input  logic sigFromSrams_bore_51_ram_bp_clken,
    input  logic sigFromSrams_bore_51_ram_aux_clk,
    input  logic sigFromSrams_bore_51_ram_aux_ckbp,
    input  logic sigFromSrams_bore_51_ram_mcp_hold,
    input  logic sigFromSrams_bore_51_cgen,
    input  logic sigFromSrams_bore_52_ram_hold,
    input  logic sigFromSrams_bore_52_ram_bypass,
    input  logic sigFromSrams_bore_52_ram_bp_clken,
    input  logic sigFromSrams_bore_52_ram_aux_clk,
    input  logic sigFromSrams_bore_52_ram_aux_ckbp,
    input  logic sigFromSrams_bore_52_ram_mcp_hold,
    input  logic sigFromSrams_bore_52_cgen,
    input  logic sigFromSrams_bore_53_ram_hold,
    input  logic sigFromSrams_bore_53_ram_bypass,
    input  logic sigFromSrams_bore_53_ram_bp_clken,
    input  logic sigFromSrams_bore_53_ram_aux_clk,
    input  logic sigFromSrams_bore_53_ram_aux_ckbp,
    input  logic sigFromSrams_bore_53_ram_mcp_hold,
    input  logic sigFromSrams_bore_53_cgen,
    input  logic sigFromSrams_bore_54_ram_hold,
    input  logic sigFromSrams_bore_54_ram_bypass,
    input  logic sigFromSrams_bore_54_ram_bp_clken,
    input  logic sigFromSrams_bore_54_ram_aux_clk,
    input  logic sigFromSrams_bore_54_ram_aux_ckbp,
    input  logic sigFromSrams_bore_54_ram_mcp_hold,
    input  logic sigFromSrams_bore_54_cgen,
    input  logic sigFromSrams_bore_55_ram_hold,
    input  logic sigFromSrams_bore_55_ram_bypass,
    input  logic sigFromSrams_bore_55_ram_bp_clken,
    input  logic sigFromSrams_bore_55_ram_aux_clk,
    input  logic sigFromSrams_bore_55_ram_aux_ckbp,
    input  logic sigFromSrams_bore_55_ram_mcp_hold,
    input  logic sigFromSrams_bore_55_cgen,
    input  logic sigFromSrams_bore_56_ram_hold,
    input  logic sigFromSrams_bore_56_ram_bypass,
    input  logic sigFromSrams_bore_56_ram_bp_clken,
    input  logic sigFromSrams_bore_56_ram_aux_clk,
    input  logic sigFromSrams_bore_56_ram_aux_ckbp,
    input  logic sigFromSrams_bore_56_ram_mcp_hold,
    input  logic sigFromSrams_bore_56_cgen,
    input  logic sigFromSrams_bore_57_ram_hold,
    input  logic sigFromSrams_bore_57_ram_bypass,
    input  logic sigFromSrams_bore_57_ram_bp_clken,
    input  logic sigFromSrams_bore_57_ram_aux_clk,
    input  logic sigFromSrams_bore_57_ram_aux_ckbp,
    input  logic sigFromSrams_bore_57_ram_mcp_hold,
    input  logic sigFromSrams_bore_57_cgen,
    input  logic sigFromSrams_bore_58_ram_hold,
    input  logic sigFromSrams_bore_58_ram_bypass,
    input  logic sigFromSrams_bore_58_ram_bp_clken,
    input  logic sigFromSrams_bore_58_ram_aux_clk,
    input  logic sigFromSrams_bore_58_ram_aux_ckbp,
    input  logic sigFromSrams_bore_58_ram_mcp_hold,
    input  logic sigFromSrams_bore_58_cgen,
    input  logic sigFromSrams_bore_59_ram_hold,
    input  logic sigFromSrams_bore_59_ram_bypass,
    input  logic sigFromSrams_bore_59_ram_bp_clken,
    input  logic sigFromSrams_bore_59_ram_aux_clk,
    input  logic sigFromSrams_bore_59_ram_aux_ckbp,
    input  logic sigFromSrams_bore_59_ram_mcp_hold,
    input  logic sigFromSrams_bore_59_cgen,
    input  logic sigFromSrams_bore_60_ram_hold,
    input  logic sigFromSrams_bore_60_ram_bypass,
    input  logic sigFromSrams_bore_60_ram_bp_clken,
    input  logic sigFromSrams_bore_60_ram_aux_clk,
    input  logic sigFromSrams_bore_60_ram_aux_ckbp,
    input  logic sigFromSrams_bore_60_ram_mcp_hold,
    input  logic sigFromSrams_bore_60_cgen,
    input  logic sigFromSrams_bore_61_ram_hold,
    input  logic sigFromSrams_bore_61_ram_bypass,
    input  logic sigFromSrams_bore_61_ram_bp_clken,
    input  logic sigFromSrams_bore_61_ram_aux_clk,
    input  logic sigFromSrams_bore_61_ram_aux_ckbp,
    input  logic sigFromSrams_bore_61_ram_mcp_hold,
    input  logic sigFromSrams_bore_61_cgen,
    input  logic sigFromSrams_bore_62_ram_hold,
    input  logic sigFromSrams_bore_62_ram_bypass,
    input  logic sigFromSrams_bore_62_ram_bp_clken,
    input  logic sigFromSrams_bore_62_ram_aux_clk,
    input  logic sigFromSrams_bore_62_ram_aux_ckbp,
    input  logic sigFromSrams_bore_62_ram_mcp_hold,
    input  logic sigFromSrams_bore_62_cgen,
    input  logic sigFromSrams_bore_63_ram_hold,
    input  logic sigFromSrams_bore_63_ram_bypass,
    input  logic sigFromSrams_bore_63_ram_bp_clken,
    input  logic sigFromSrams_bore_63_ram_aux_clk,
    input  logic sigFromSrams_bore_63_ram_aux_ckbp,
    input  logic sigFromSrams_bore_63_ram_mcp_hold,
    input  logic sigFromSrams_bore_63_cgen,
    input  logic sigFromSrams_bore_64_ram_hold,
    input  logic sigFromSrams_bore_64_ram_bypass,
    input  logic sigFromSrams_bore_64_ram_bp_clken,
    input  logic sigFromSrams_bore_64_ram_aux_clk,
    input  logic sigFromSrams_bore_64_ram_aux_ckbp,
    input  logic sigFromSrams_bore_64_ram_mcp_hold,
    input  logic sigFromSrams_bore_64_cgen,
    input  logic sigFromSrams_bore_65_ram_hold,
    input  logic sigFromSrams_bore_65_ram_bypass,
    input  logic sigFromSrams_bore_65_ram_bp_clken,
    input  logic sigFromSrams_bore_65_ram_aux_clk,
    input  logic sigFromSrams_bore_65_ram_aux_ckbp,
    input  logic sigFromSrams_bore_65_ram_mcp_hold,
    input  logic sigFromSrams_bore_65_cgen,
    input  logic sigFromSrams_bore_66_ram_hold,
    input  logic sigFromSrams_bore_66_ram_bypass,
    input  logic sigFromSrams_bore_66_ram_bp_clken,
    input  logic sigFromSrams_bore_66_ram_aux_clk,
    input  logic sigFromSrams_bore_66_ram_aux_ckbp,
    input  logic sigFromSrams_bore_66_ram_mcp_hold,
    input  logic sigFromSrams_bore_66_cgen,
    input  logic sigFromSrams_bore_67_ram_hold,
    input  logic sigFromSrams_bore_67_ram_bypass,
    input  logic sigFromSrams_bore_67_ram_bp_clken,
    input  logic sigFromSrams_bore_67_ram_aux_clk,
    input  logic sigFromSrams_bore_67_ram_aux_ckbp,
    input  logic sigFromSrams_bore_67_ram_mcp_hold,
    input  logic sigFromSrams_bore_67_cgen,
    input  logic sigFromSrams_bore_68_ram_hold,
    input  logic sigFromSrams_bore_68_ram_bypass,
    input  logic sigFromSrams_bore_68_ram_bp_clken,
    input  logic sigFromSrams_bore_68_ram_aux_clk,
    input  logic sigFromSrams_bore_68_ram_aux_ckbp,
    input  logic sigFromSrams_bore_68_ram_mcp_hold,
    input  logic sigFromSrams_bore_68_cgen,
    input  logic sigFromSrams_bore_69_ram_hold,
    input  logic sigFromSrams_bore_69_ram_bypass,
    input  logic sigFromSrams_bore_69_ram_bp_clken,
    input  logic sigFromSrams_bore_69_ram_aux_clk,
    input  logic sigFromSrams_bore_69_ram_aux_ckbp,
    input  logic sigFromSrams_bore_69_ram_mcp_hold,
    input  logic sigFromSrams_bore_69_cgen,
    input  logic sigFromSrams_bore_70_ram_hold,
    input  logic sigFromSrams_bore_70_ram_bypass,
    input  logic sigFromSrams_bore_70_ram_bp_clken,
    input  logic sigFromSrams_bore_70_ram_aux_clk,
    input  logic sigFromSrams_bore_70_ram_aux_ckbp,
    input  logic sigFromSrams_bore_70_ram_mcp_hold,
    input  logic sigFromSrams_bore_70_cgen,
    input  logic sigFromSrams_bore_71_ram_hold,
    input  logic sigFromSrams_bore_71_ram_bypass,
    input  logic sigFromSrams_bore_71_ram_bp_clken,
    input  logic sigFromSrams_bore_71_ram_aux_clk,
    input  logic sigFromSrams_bore_71_ram_aux_ckbp,
    input  logic sigFromSrams_bore_71_ram_mcp_hold,
    input  logic sigFromSrams_bore_71_cgen,
    input  logic sigFromSrams_bore_72_ram_hold,
    input  logic sigFromSrams_bore_72_ram_bypass,
    input  logic sigFromSrams_bore_72_ram_bp_clken,
    input  logic sigFromSrams_bore_72_ram_aux_clk,
    input  logic sigFromSrams_bore_72_ram_aux_ckbp,
    input  logic sigFromSrams_bore_72_ram_mcp_hold,
    input  logic sigFromSrams_bore_72_cgen,
    input  logic sigFromSrams_bore_73_ram_hold,
    input  logic sigFromSrams_bore_73_ram_bypass,
    input  logic sigFromSrams_bore_73_ram_bp_clken,
    input  logic sigFromSrams_bore_73_ram_aux_clk,
    input  logic sigFromSrams_bore_73_ram_aux_ckbp,
    input  logic sigFromSrams_bore_73_ram_mcp_hold,
    input  logic sigFromSrams_bore_73_cgen,
    input  logic sigFromSrams_bore_74_ram_hold,
    input  logic sigFromSrams_bore_74_ram_bypass,
    input  logic sigFromSrams_bore_74_ram_bp_clken,
    input  logic sigFromSrams_bore_74_ram_aux_clk,
    input  logic sigFromSrams_bore_74_ram_aux_ckbp,
    input  logic sigFromSrams_bore_74_ram_mcp_hold,
    input  logic sigFromSrams_bore_74_cgen,
    input  logic sigFromSrams_bore_75_ram_hold,
    input  logic sigFromSrams_bore_75_ram_bypass,
    input  logic sigFromSrams_bore_75_ram_bp_clken,
    input  logic sigFromSrams_bore_75_ram_aux_clk,
    input  logic sigFromSrams_bore_75_ram_aux_ckbp,
    input  logic sigFromSrams_bore_75_ram_mcp_hold,
    input  logic sigFromSrams_bore_75_cgen,
    input  logic sigFromSrams_bore_76_ram_hold,
    input  logic sigFromSrams_bore_76_ram_bypass,
    input  logic sigFromSrams_bore_76_ram_bp_clken,
    input  logic sigFromSrams_bore_76_ram_aux_clk,
    input  logic sigFromSrams_bore_76_ram_aux_ckbp,
    input  logic sigFromSrams_bore_76_ram_mcp_hold,
    input  logic sigFromSrams_bore_76_cgen,
    input  logic sigFromSrams_bore_77_ram_hold,
    input  logic sigFromSrams_bore_77_ram_bypass,
    input  logic sigFromSrams_bore_77_ram_bp_clken,
    input  logic sigFromSrams_bore_77_ram_aux_clk,
    input  logic sigFromSrams_bore_77_ram_aux_ckbp,
    input  logic sigFromSrams_bore_77_ram_mcp_hold,
    input  logic sigFromSrams_bore_77_cgen,
    input  logic sigFromSrams_bore_78_ram_hold,
    input  logic sigFromSrams_bore_78_ram_bypass,
    input  logic sigFromSrams_bore_78_ram_bp_clken,
    input  logic sigFromSrams_bore_78_ram_aux_clk,
    input  logic sigFromSrams_bore_78_ram_aux_ckbp,
    input  logic sigFromSrams_bore_78_ram_mcp_hold,
    input  logic sigFromSrams_bore_78_cgen,
    input  logic sigFromSrams_bore_79_ram_hold,
    input  logic sigFromSrams_bore_79_ram_bypass,
    input  logic sigFromSrams_bore_79_ram_bp_clken,
    input  logic sigFromSrams_bore_79_ram_aux_clk,
    input  logic sigFromSrams_bore_79_ram_aux_ckbp,
    input  logic sigFromSrams_bore_79_ram_mcp_hold,
    input  logic sigFromSrams_bore_79_cgen,
    input  logic sigFromSrams_bore_80_ram_hold,
    input  logic sigFromSrams_bore_80_ram_bypass,
    input  logic sigFromSrams_bore_80_ram_bp_clken,
    input  logic sigFromSrams_bore_80_ram_aux_clk,
    input  logic sigFromSrams_bore_80_ram_aux_ckbp,
    input  logic sigFromSrams_bore_80_ram_mcp_hold,
    input  logic sigFromSrams_bore_80_cgen,
    input  logic sigFromSrams_bore_81_ram_hold,
    input  logic sigFromSrams_bore_81_ram_bypass,
    input  logic sigFromSrams_bore_81_ram_bp_clken,
    input  logic sigFromSrams_bore_81_ram_aux_clk,
    input  logic sigFromSrams_bore_81_ram_aux_ckbp,
    input  logic sigFromSrams_bore_81_ram_mcp_hold,
    input  logic sigFromSrams_bore_81_cgen,
    input  logic sigFromSrams_bore_82_ram_hold,
    input  logic sigFromSrams_bore_82_ram_bypass,
    input  logic sigFromSrams_bore_82_ram_bp_clken,
    input  logic sigFromSrams_bore_82_ram_aux_clk,
    input  logic sigFromSrams_bore_82_ram_aux_ckbp,
    input  logic sigFromSrams_bore_82_ram_mcp_hold,
    input  logic sigFromSrams_bore_82_cgen,
    input  logic sigFromSrams_bore_83_ram_hold,
    input  logic sigFromSrams_bore_83_ram_bypass,
    input  logic sigFromSrams_bore_83_ram_bp_clken,
    input  logic sigFromSrams_bore_83_ram_aux_clk,
    input  logic sigFromSrams_bore_83_ram_aux_ckbp,
    input  logic sigFromSrams_bore_83_ram_mcp_hold,
    input  logic sigFromSrams_bore_83_cgen,
    input  logic sigFromSrams_bore_84_ram_hold,
    input  logic sigFromSrams_bore_84_ram_bypass,
    input  logic sigFromSrams_bore_84_ram_bp_clken,
    input  logic sigFromSrams_bore_84_ram_aux_clk,
    input  logic sigFromSrams_bore_84_ram_aux_ckbp,
    input  logic sigFromSrams_bore_84_ram_mcp_hold,
    input  logic sigFromSrams_bore_84_cgen,
    input  logic sigFromSrams_bore_85_ram_hold,
    input  logic sigFromSrams_bore_85_ram_bypass,
    input  logic sigFromSrams_bore_85_ram_bp_clken,
    input  logic sigFromSrams_bore_85_ram_aux_clk,
    input  logic sigFromSrams_bore_85_ram_aux_ckbp,
    input  logic sigFromSrams_bore_85_ram_mcp_hold,
    input  logic sigFromSrams_bore_85_cgen,
    input  logic sigFromSrams_bore_86_ram_hold,
    input  logic sigFromSrams_bore_86_ram_bypass,
    input  logic sigFromSrams_bore_86_ram_bp_clken,
    input  logic sigFromSrams_bore_86_ram_aux_clk,
    input  logic sigFromSrams_bore_86_ram_aux_ckbp,
    input  logic sigFromSrams_bore_86_ram_mcp_hold,
    input  logic sigFromSrams_bore_86_cgen,
    input  logic sigFromSrams_bore_87_ram_hold,
    input  logic sigFromSrams_bore_87_ram_bypass,
    input  logic sigFromSrams_bore_87_ram_bp_clken,
    input  logic sigFromSrams_bore_87_ram_aux_clk,
    input  logic sigFromSrams_bore_87_ram_aux_ckbp,
    input  logic sigFromSrams_bore_87_ram_mcp_hold,
    input  logic sigFromSrams_bore_87_cgen,
    input  logic sigFromSrams_bore_88_ram_hold,
    input  logic sigFromSrams_bore_88_ram_bypass,
    input  logic sigFromSrams_bore_88_ram_bp_clken,
    input  logic sigFromSrams_bore_88_ram_aux_clk,
    input  logic sigFromSrams_bore_88_ram_aux_ckbp,
    input  logic sigFromSrams_bore_88_ram_mcp_hold,
    input  logic sigFromSrams_bore_88_cgen,
    input  logic sigFromSrams_bore_89_ram_hold,
    input  logic sigFromSrams_bore_89_ram_bypass,
    input  logic sigFromSrams_bore_89_ram_bp_clken,
    input  logic sigFromSrams_bore_89_ram_aux_clk,
    input  logic sigFromSrams_bore_89_ram_aux_ckbp,
    input  logic sigFromSrams_bore_89_ram_mcp_hold,
    input  logic sigFromSrams_bore_89_cgen,
    input  logic sigFromSrams_bore_90_ram_hold,
    input  logic sigFromSrams_bore_90_ram_bypass,
    input  logic sigFromSrams_bore_90_ram_bp_clken,
    input  logic sigFromSrams_bore_90_ram_aux_clk,
    input  logic sigFromSrams_bore_90_ram_aux_ckbp,
    input  logic sigFromSrams_bore_90_ram_mcp_hold,
    input  logic sigFromSrams_bore_90_cgen,
    input  logic sigFromSrams_bore_91_ram_hold,
    input  logic sigFromSrams_bore_91_ram_bypass,
    input  logic sigFromSrams_bore_91_ram_bp_clken,
    input  logic sigFromSrams_bore_91_ram_aux_clk,
    input  logic sigFromSrams_bore_91_ram_aux_ckbp,
    input  logic sigFromSrams_bore_91_ram_mcp_hold,
    input  logic sigFromSrams_bore_91_cgen,
    input  logic sigFromSrams_bore_92_ram_hold,
    input  logic sigFromSrams_bore_92_ram_bypass,
    input  logic sigFromSrams_bore_92_ram_bp_clken,
    input  logic sigFromSrams_bore_92_ram_aux_clk,
    input  logic sigFromSrams_bore_92_ram_aux_ckbp,
    input  logic sigFromSrams_bore_92_ram_mcp_hold,
    input  logic sigFromSrams_bore_92_cgen,
    input  logic sigFromSrams_bore_93_ram_hold,
    input  logic sigFromSrams_bore_93_ram_bypass,
    input  logic sigFromSrams_bore_93_ram_bp_clken,
    input  logic sigFromSrams_bore_93_ram_aux_clk,
    input  logic sigFromSrams_bore_93_ram_aux_ckbp,
    input  logic sigFromSrams_bore_93_ram_mcp_hold,
    input  logic sigFromSrams_bore_93_cgen,
    input  logic sigFromSrams_bore_94_ram_hold,
    input  logic sigFromSrams_bore_94_ram_bypass,
    input  logic sigFromSrams_bore_94_ram_bp_clken,
    input  logic sigFromSrams_bore_94_ram_aux_clk,
    input  logic sigFromSrams_bore_94_ram_aux_ckbp,
    input  logic sigFromSrams_bore_94_ram_mcp_hold,
    input  logic sigFromSrams_bore_94_cgen,
    input  logic sigFromSrams_bore_95_ram_hold,
    input  logic sigFromSrams_bore_95_ram_bypass,
    input  logic sigFromSrams_bore_95_ram_bp_clken,
    input  logic sigFromSrams_bore_95_ram_aux_clk,
    input  logic sigFromSrams_bore_95_ram_aux_ckbp,
    input  logic sigFromSrams_bore_95_ram_mcp_hold,
    input  logic sigFromSrams_bore_95_cgen,
    input  logic sigFromSrams_bore_96_ram_hold,
    input  logic sigFromSrams_bore_96_ram_bypass,
    input  logic sigFromSrams_bore_96_ram_bp_clken,
    input  logic sigFromSrams_bore_96_ram_aux_clk,
    input  logic sigFromSrams_bore_96_ram_aux_ckbp,
    input  logic sigFromSrams_bore_96_ram_mcp_hold,
    input  logic sigFromSrams_bore_96_cgen,
    input  logic sigFromSrams_bore_97_ram_hold,
    input  logic sigFromSrams_bore_97_ram_bypass,
    input  logic sigFromSrams_bore_97_ram_bp_clken,
    input  logic sigFromSrams_bore_97_ram_aux_clk,
    input  logic sigFromSrams_bore_97_ram_aux_ckbp,
    input  logic sigFromSrams_bore_97_ram_mcp_hold,
    input  logic sigFromSrams_bore_97_cgen,
    input  logic sigFromSrams_bore_98_ram_hold,
    input  logic sigFromSrams_bore_98_ram_bypass,
    input  logic sigFromSrams_bore_98_ram_bp_clken,
    input  logic sigFromSrams_bore_98_ram_aux_clk,
    input  logic sigFromSrams_bore_98_ram_aux_ckbp,
    input  logic sigFromSrams_bore_98_ram_mcp_hold,
    input  logic sigFromSrams_bore_98_cgen,
    input  logic sigFromSrams_bore_99_ram_hold,
    input  logic sigFromSrams_bore_99_ram_bypass,
    input  logic sigFromSrams_bore_99_ram_bp_clken,
    input  logic sigFromSrams_bore_99_ram_aux_clk,
    input  logic sigFromSrams_bore_99_ram_aux_ckbp,
    input  logic sigFromSrams_bore_99_ram_mcp_hold,
    input  logic sigFromSrams_bore_99_cgen,
    input  logic sigFromSrams_bore_100_ram_hold,
    input  logic sigFromSrams_bore_100_ram_bypass,
    input  logic sigFromSrams_bore_100_ram_bp_clken,
    input  logic sigFromSrams_bore_100_ram_aux_clk,
    input  logic sigFromSrams_bore_100_ram_aux_ckbp,
    input  logic sigFromSrams_bore_100_ram_mcp_hold,
    input  logic sigFromSrams_bore_100_cgen,
    input  logic sigFromSrams_bore_101_ram_hold,
    input  logic sigFromSrams_bore_101_ram_bypass,
    input  logic sigFromSrams_bore_101_ram_bp_clken,
    input  logic sigFromSrams_bore_101_ram_aux_clk,
    input  logic sigFromSrams_bore_101_ram_aux_ckbp,
    input  logic sigFromSrams_bore_101_ram_mcp_hold,
    input  logic sigFromSrams_bore_101_cgen,
    input  logic sigFromSrams_bore_102_ram_hold,
    input  logic sigFromSrams_bore_102_ram_bypass,
    input  logic sigFromSrams_bore_102_ram_bp_clken,
    input  logic sigFromSrams_bore_102_ram_aux_clk,
    input  logic sigFromSrams_bore_102_ram_aux_ckbp,
    input  logic sigFromSrams_bore_102_ram_mcp_hold,
    input  logic sigFromSrams_bore_102_cgen,
    input  logic sigFromSrams_bore_103_ram_hold,
    input  logic sigFromSrams_bore_103_ram_bypass,
    input  logic sigFromSrams_bore_103_ram_bp_clken,
    input  logic sigFromSrams_bore_103_ram_aux_clk,
    input  logic sigFromSrams_bore_103_ram_aux_ckbp,
    input  logic sigFromSrams_bore_103_ram_mcp_hold,
    input  logic sigFromSrams_bore_103_cgen,
    input  logic sigFromSrams_bore_104_ram_hold,
    input  logic sigFromSrams_bore_104_ram_bypass,
    input  logic sigFromSrams_bore_104_ram_bp_clken,
    input  logic sigFromSrams_bore_104_ram_aux_clk,
    input  logic sigFromSrams_bore_104_ram_aux_ckbp,
    input  logic sigFromSrams_bore_104_ram_mcp_hold,
    input  logic sigFromSrams_bore_104_cgen,
    input  logic sigFromSrams_bore_105_ram_hold,
    input  logic sigFromSrams_bore_105_ram_bypass,
    input  logic sigFromSrams_bore_105_ram_bp_clken,
    input  logic sigFromSrams_bore_105_ram_aux_clk,
    input  logic sigFromSrams_bore_105_ram_aux_ckbp,
    input  logic sigFromSrams_bore_105_ram_mcp_hold,
    input  logic sigFromSrams_bore_105_cgen,
    input  logic sigFromSrams_bore_106_ram_hold,
    input  logic sigFromSrams_bore_106_ram_bypass,
    input  logic sigFromSrams_bore_106_ram_bp_clken,
    input  logic sigFromSrams_bore_106_ram_aux_clk,
    input  logic sigFromSrams_bore_106_ram_aux_ckbp,
    input  logic sigFromSrams_bore_106_ram_mcp_hold,
    input  logic sigFromSrams_bore_106_cgen,
    input  logic sigFromSrams_bore_107_ram_hold,
    input  logic sigFromSrams_bore_107_ram_bypass,
    input  logic sigFromSrams_bore_107_ram_bp_clken,
    input  logic sigFromSrams_bore_107_ram_aux_clk,
    input  logic sigFromSrams_bore_107_ram_aux_ckbp,
    input  logic sigFromSrams_bore_107_ram_mcp_hold,
    input  logic sigFromSrams_bore_107_cgen,
    input  logic sigFromSrams_bore_108_ram_hold,
    input  logic sigFromSrams_bore_108_ram_bypass,
    input  logic sigFromSrams_bore_108_ram_bp_clken,
    input  logic sigFromSrams_bore_108_ram_aux_clk,
    input  logic sigFromSrams_bore_108_ram_aux_ckbp,
    input  logic sigFromSrams_bore_108_ram_mcp_hold,
    input  logic sigFromSrams_bore_108_cgen,
    input  logic sigFromSrams_bore_109_ram_hold,
    input  logic sigFromSrams_bore_109_ram_bypass,
    input  logic sigFromSrams_bore_109_ram_bp_clken,
    input  logic sigFromSrams_bore_109_ram_aux_clk,
    input  logic sigFromSrams_bore_109_ram_aux_ckbp,
    input  logic sigFromSrams_bore_109_ram_mcp_hold,
    input  logic sigFromSrams_bore_109_cgen,
    input  logic sigFromSrams_bore_110_ram_hold,
    input  logic sigFromSrams_bore_110_ram_bypass,
    input  logic sigFromSrams_bore_110_ram_bp_clken,
    input  logic sigFromSrams_bore_110_ram_aux_clk,
    input  logic sigFromSrams_bore_110_ram_aux_ckbp,
    input  logic sigFromSrams_bore_110_ram_mcp_hold,
    input  logic sigFromSrams_bore_110_cgen,
    input  logic sigFromSrams_bore_111_ram_hold,
    input  logic sigFromSrams_bore_111_ram_bypass,
    input  logic sigFromSrams_bore_111_ram_bp_clken,
    input  logic sigFromSrams_bore_111_ram_aux_clk,
    input  logic sigFromSrams_bore_111_ram_aux_ckbp,
    input  logic sigFromSrams_bore_111_ram_mcp_hold,
    input  logic sigFromSrams_bore_111_cgen,
    input  logic sigFromSrams_bore_112_ram_hold,
    input  logic sigFromSrams_bore_112_ram_bypass,
    input  logic sigFromSrams_bore_112_ram_bp_clken,
    input  logic sigFromSrams_bore_112_ram_aux_clk,
    input  logic sigFromSrams_bore_112_ram_aux_ckbp,
    input  logic sigFromSrams_bore_112_ram_mcp_hold,
    input  logic sigFromSrams_bore_112_cgen,
    input  logic sigFromSrams_bore_113_ram_hold,
    input  logic sigFromSrams_bore_113_ram_bypass,
    input  logic sigFromSrams_bore_113_ram_bp_clken,
    input  logic sigFromSrams_bore_113_ram_aux_clk,
    input  logic sigFromSrams_bore_113_ram_aux_ckbp,
    input  logic sigFromSrams_bore_113_ram_mcp_hold,
    input  logic sigFromSrams_bore_113_cgen,
    input  logic sigFromSrams_bore_114_ram_hold,
    input  logic sigFromSrams_bore_114_ram_bypass,
    input  logic sigFromSrams_bore_114_ram_bp_clken,
    input  logic sigFromSrams_bore_114_ram_aux_clk,
    input  logic sigFromSrams_bore_114_ram_aux_ckbp,
    input  logic sigFromSrams_bore_114_ram_mcp_hold,
    input  logic sigFromSrams_bore_114_cgen,
    input  logic sigFromSrams_bore_115_ram_hold,
    input  logic sigFromSrams_bore_115_ram_bypass,
    input  logic sigFromSrams_bore_115_ram_bp_clken,
    input  logic sigFromSrams_bore_115_ram_aux_clk,
    input  logic sigFromSrams_bore_115_ram_aux_ckbp,
    input  logic sigFromSrams_bore_115_ram_mcp_hold,
    input  logic sigFromSrams_bore_115_cgen,
    input  logic sigFromSrams_bore_116_ram_hold,
    input  logic sigFromSrams_bore_116_ram_bypass,
    input  logic sigFromSrams_bore_116_ram_bp_clken,
    input  logic sigFromSrams_bore_116_ram_aux_clk,
    input  logic sigFromSrams_bore_116_ram_aux_ckbp,
    input  logic sigFromSrams_bore_116_ram_mcp_hold,
    input  logic sigFromSrams_bore_116_cgen,
    input  logic sigFromSrams_bore_117_ram_hold,
    input  logic sigFromSrams_bore_117_ram_bypass,
    input  logic sigFromSrams_bore_117_ram_bp_clken,
    input  logic sigFromSrams_bore_117_ram_aux_clk,
    input  logic sigFromSrams_bore_117_ram_aux_ckbp,
    input  logic sigFromSrams_bore_117_ram_mcp_hold,
    input  logic sigFromSrams_bore_117_cgen,
    input  logic sigFromSrams_bore_118_ram_hold,
    input  logic sigFromSrams_bore_118_ram_bypass,
    input  logic sigFromSrams_bore_118_ram_bp_clken,
    input  logic sigFromSrams_bore_118_ram_aux_clk,
    input  logic sigFromSrams_bore_118_ram_aux_ckbp,
    input  logic sigFromSrams_bore_118_ram_mcp_hold,
    input  logic sigFromSrams_bore_118_cgen,
    input  logic sigFromSrams_bore_119_ram_hold,
    input  logic sigFromSrams_bore_119_ram_bypass,
    input  logic sigFromSrams_bore_119_ram_bp_clken,
    input  logic sigFromSrams_bore_119_ram_aux_clk,
    input  logic sigFromSrams_bore_119_ram_aux_ckbp,
    input  logic sigFromSrams_bore_119_ram_mcp_hold,
    input  logic sigFromSrams_bore_119_cgen,
    input  logic sigFromSrams_bore_120_ram_hold,
    input  logic sigFromSrams_bore_120_ram_bypass,
    input  logic sigFromSrams_bore_120_ram_bp_clken,
    input  logic sigFromSrams_bore_120_ram_aux_clk,
    input  logic sigFromSrams_bore_120_ram_aux_ckbp,
    input  logic sigFromSrams_bore_120_ram_mcp_hold,
    input  logic sigFromSrams_bore_120_cgen,
    input  logic sigFromSrams_bore_121_ram_hold,
    input  logic sigFromSrams_bore_121_ram_bypass,
    input  logic sigFromSrams_bore_121_ram_bp_clken,
    input  logic sigFromSrams_bore_121_ram_aux_clk,
    input  logic sigFromSrams_bore_121_ram_aux_ckbp,
    input  logic sigFromSrams_bore_121_ram_mcp_hold,
    input  logic sigFromSrams_bore_121_cgen,
    input  logic sigFromSrams_bore_122_ram_hold,
    input  logic sigFromSrams_bore_122_ram_bypass,
    input  logic sigFromSrams_bore_122_ram_bp_clken,
    input  logic sigFromSrams_bore_122_ram_aux_clk,
    input  logic sigFromSrams_bore_122_ram_aux_ckbp,
    input  logic sigFromSrams_bore_122_ram_mcp_hold,
    input  logic sigFromSrams_bore_122_cgen,
    input  logic sigFromSrams_bore_123_ram_hold,
    input  logic sigFromSrams_bore_123_ram_bypass,
    input  logic sigFromSrams_bore_123_ram_bp_clken,
    input  logic sigFromSrams_bore_123_ram_aux_clk,
    input  logic sigFromSrams_bore_123_ram_aux_ckbp,
    input  logic sigFromSrams_bore_123_ram_mcp_hold,
    input  logic sigFromSrams_bore_123_cgen,
    input  logic sigFromSrams_bore_124_ram_hold,
    input  logic sigFromSrams_bore_124_ram_bypass,
    input  logic sigFromSrams_bore_124_ram_bp_clken,
    input  logic sigFromSrams_bore_124_ram_aux_clk,
    input  logic sigFromSrams_bore_124_ram_aux_ckbp,
    input  logic sigFromSrams_bore_124_ram_mcp_hold,
    input  logic sigFromSrams_bore_124_cgen,
    input  logic sigFromSrams_bore_125_ram_hold,
    input  logic sigFromSrams_bore_125_ram_bypass,
    input  logic sigFromSrams_bore_125_ram_bp_clken,
    input  logic sigFromSrams_bore_125_ram_aux_clk,
    input  logic sigFromSrams_bore_125_ram_aux_ckbp,
    input  logic sigFromSrams_bore_125_ram_mcp_hold,
    input  logic sigFromSrams_bore_125_cgen,
    input  logic sigFromSrams_bore_126_ram_hold,
    input  logic sigFromSrams_bore_126_ram_bypass,
    input  logic sigFromSrams_bore_126_ram_bp_clken,
    input  logic sigFromSrams_bore_126_ram_aux_clk,
    input  logic sigFromSrams_bore_126_ram_aux_ckbp,
    input  logic sigFromSrams_bore_126_ram_mcp_hold,
    input  logic sigFromSrams_bore_126_cgen,
    input  logic sigFromSrams_bore_127_ram_hold,
    input  logic sigFromSrams_bore_127_ram_bypass,
    input  logic sigFromSrams_bore_127_ram_bp_clken,
    input  logic sigFromSrams_bore_127_ram_aux_clk,
    input  logic sigFromSrams_bore_127_ram_aux_ckbp,
    input  logic sigFromSrams_bore_127_ram_mcp_hold,
    input  logic sigFromSrams_bore_127_cgen,
    input  logic sigFromSrams_bore_128_ram_hold,
    input  logic sigFromSrams_bore_128_ram_bypass,
    input  logic sigFromSrams_bore_128_ram_bp_clken,
    input  logic sigFromSrams_bore_128_ram_aux_clk,
    input  logic sigFromSrams_bore_128_ram_aux_ckbp,
    input  logic sigFromSrams_bore_128_ram_mcp_hold,
    input  logic sigFromSrams_bore_128_cgen,
    input  logic sigFromSrams_bore_129_ram_hold,
    input  logic sigFromSrams_bore_129_ram_bypass,
    input  logic sigFromSrams_bore_129_ram_bp_clken,
    input  logic sigFromSrams_bore_129_ram_aux_clk,
    input  logic sigFromSrams_bore_129_ram_aux_ckbp,
    input  logic sigFromSrams_bore_129_ram_mcp_hold,
    input  logic sigFromSrams_bore_129_cgen,
    input  logic sigFromSrams_bore_130_ram_hold,
    input  logic sigFromSrams_bore_130_ram_bypass,
    input  logic sigFromSrams_bore_130_ram_bp_clken,
    input  logic sigFromSrams_bore_130_ram_aux_clk,
    input  logic sigFromSrams_bore_130_ram_aux_ckbp,
    input  logic sigFromSrams_bore_130_ram_mcp_hold,
    input  logic sigFromSrams_bore_130_cgen,
    input  logic sigFromSrams_bore_131_ram_hold,
    input  logic sigFromSrams_bore_131_ram_bypass,
    input  logic sigFromSrams_bore_131_ram_bp_clken,
    input  logic sigFromSrams_bore_131_ram_aux_clk,
    input  logic sigFromSrams_bore_131_ram_aux_ckbp,
    input  logic sigFromSrams_bore_131_ram_mcp_hold,
    input  logic sigFromSrams_bore_131_cgen,
    input  logic sigFromSrams_bore_132_ram_hold,
    input  logic sigFromSrams_bore_132_ram_bypass,
    input  logic sigFromSrams_bore_132_ram_bp_clken,
    input  logic sigFromSrams_bore_132_ram_aux_clk,
    input  logic sigFromSrams_bore_132_ram_aux_ckbp,
    input  logic sigFromSrams_bore_132_ram_mcp_hold,
    input  logic sigFromSrams_bore_132_cgen,
    input  logic sigFromSrams_bore_133_ram_hold,
    input  logic sigFromSrams_bore_133_ram_bypass,
    input  logic sigFromSrams_bore_133_ram_bp_clken,
    input  logic sigFromSrams_bore_133_ram_aux_clk,
    input  logic sigFromSrams_bore_133_ram_aux_ckbp,
    input  logic sigFromSrams_bore_133_ram_mcp_hold,
    input  logic sigFromSrams_bore_133_cgen,
    input  logic sigFromSrams_bore_134_ram_hold,
    input  logic sigFromSrams_bore_134_ram_bypass,
    input  logic sigFromSrams_bore_134_ram_bp_clken,
    input  logic sigFromSrams_bore_134_ram_aux_clk,
    input  logic sigFromSrams_bore_134_ram_aux_ckbp,
    input  logic sigFromSrams_bore_134_ram_mcp_hold,
    input  logic sigFromSrams_bore_134_cgen,
    input  logic sigFromSrams_bore_135_ram_hold,
    input  logic sigFromSrams_bore_135_ram_bypass,
    input  logic sigFromSrams_bore_135_ram_bp_clken,
    input  logic sigFromSrams_bore_135_ram_aux_clk,
    input  logic sigFromSrams_bore_135_ram_aux_ckbp,
    input  logic sigFromSrams_bore_135_ram_mcp_hold,
    input  logic sigFromSrams_bore_135_cgen,
    input  logic sigFromSrams_bore_136_ram_hold,
    input  logic sigFromSrams_bore_136_ram_bypass,
    input  logic sigFromSrams_bore_136_ram_bp_clken,
    input  logic sigFromSrams_bore_136_ram_aux_clk,
    input  logic sigFromSrams_bore_136_ram_aux_ckbp,
    input  logic sigFromSrams_bore_136_ram_mcp_hold,
    input  logic sigFromSrams_bore_136_cgen,
    input  logic sigFromSrams_bore_137_ram_hold,
    input  logic sigFromSrams_bore_137_ram_bypass,
    input  logic sigFromSrams_bore_137_ram_bp_clken,
    input  logic sigFromSrams_bore_137_ram_aux_clk,
    input  logic sigFromSrams_bore_137_ram_aux_ckbp,
    input  logic sigFromSrams_bore_137_ram_mcp_hold,
    input  logic sigFromSrams_bore_137_cgen,
    input  logic sigFromSrams_bore_138_ram_hold,
    input  logic sigFromSrams_bore_138_ram_bypass,
    input  logic sigFromSrams_bore_138_ram_bp_clken,
    input  logic sigFromSrams_bore_138_ram_aux_clk,
    input  logic sigFromSrams_bore_138_ram_aux_ckbp,
    input  logic sigFromSrams_bore_138_ram_mcp_hold,
    input  logic sigFromSrams_bore_138_cgen,
    input  logic sigFromSrams_bore_139_ram_hold,
    input  logic sigFromSrams_bore_139_ram_bypass,
    input  logic sigFromSrams_bore_139_ram_bp_clken,
    input  logic sigFromSrams_bore_139_ram_aux_clk,
    input  logic sigFromSrams_bore_139_ram_aux_ckbp,
    input  logic sigFromSrams_bore_139_ram_mcp_hold,
    input  logic sigFromSrams_bore_139_cgen,
    input  logic sigFromSrams_bore_140_ram_hold,
    input  logic sigFromSrams_bore_140_ram_bypass,
    input  logic sigFromSrams_bore_140_ram_bp_clken,
    input  logic sigFromSrams_bore_140_ram_aux_clk,
    input  logic sigFromSrams_bore_140_ram_aux_ckbp,
    input  logic sigFromSrams_bore_140_ram_mcp_hold,
    input  logic sigFromSrams_bore_140_cgen,
    input  logic sigFromSrams_bore_141_ram_hold,
    input  logic sigFromSrams_bore_141_ram_bypass,
    input  logic sigFromSrams_bore_141_ram_bp_clken,
    input  logic sigFromSrams_bore_141_ram_aux_clk,
    input  logic sigFromSrams_bore_141_ram_aux_ckbp,
    input  logic sigFromSrams_bore_141_ram_mcp_hold,
    input  logic sigFromSrams_bore_141_cgen,
    input  logic sigFromSrams_bore_142_ram_hold,
    input  logic sigFromSrams_bore_142_ram_bypass,
    input  logic sigFromSrams_bore_142_ram_bp_clken,
    input  logic sigFromSrams_bore_142_ram_aux_clk,
    input  logic sigFromSrams_bore_142_ram_aux_ckbp,
    input  logic sigFromSrams_bore_142_ram_mcp_hold,
    input  logic sigFromSrams_bore_142_cgen,
    input  logic sigFromSrams_bore_143_ram_hold,
    input  logic sigFromSrams_bore_143_ram_bypass,
    input  logic sigFromSrams_bore_143_ram_bp_clken,
    input  logic sigFromSrams_bore_143_ram_aux_clk,
    input  logic sigFromSrams_bore_143_ram_aux_ckbp,
    input  logic sigFromSrams_bore_143_ram_mcp_hold,
    input  logic sigFromSrams_bore_143_cgen,
    output logic io_toFtq_prediction_ready_o,
    output logic s1_fire_o,
    output logic abtb_io_stageCtrl_s0_fire_probe_o
);

    logic io_fromFtq_train_ready;
    logic io_toFtq_prediction_valid;
    logic [48:0] io_toFtq_prediction_bits_startPc_addr;
    logic [48:0] io_toFtq_prediction_bits_target_addr;
    logic io_toFtq_prediction_bits_takenCfiOffset_valid;
    logic [4:0] io_toFtq_prediction_bits_takenCfiOffset_bits;
    logic io_toFtq_prediction_bits_s3Override;
    logic io_toFtq_meta_valid;
    logic io_toFtq_meta_bits_redirectMeta_phr_phrPtr_flag;
    logic [9:0] io_toFtq_meta_bits_redirectMeta_phr_phrPtr_value;
    logic [12:0] io_toFtq_meta_bits_redirectMeta_phr_phrLowBits;
    logic [15:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_ghr;
    logic [7:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_bw;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_0;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_1;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_2;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_3;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_4;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_5;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_6;
    logic io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_7;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_0_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_1_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_2_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_3_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_4_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_5_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_6_branchType;
    logic [1:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_7_branchType;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_0;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_1;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_2;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_3;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_4;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_5;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_6;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_7;
    logic [3:0] io_toFtq_meta_bits_redirectMeta_ras_ssp;
    logic [2:0] io_toFtq_meta_bits_redirectMeta_ras_sctr;
    logic io_toFtq_meta_bits_redirectMeta_ras_tosw_flag;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_ras_tosw_value;
    logic io_toFtq_meta_bits_redirectMeta_ras_tosr_flag;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_ras_tosr_value;
    logic io_toFtq_meta_bits_redirectMeta_ras_nos_flag;
    logic [4:0] io_toFtq_meta_bits_redirectMeta_ras_nos_value;
    logic [48:0] io_toFtq_meta_bits_redirectMeta_ras_topRetAddr_addr;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_rawHit;
    logic [4:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_position;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_attribute_branchType;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_attribute_rasAction;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_counter_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_0_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_0_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_1_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_1_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_2_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_2_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_3_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_3_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_4_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_4_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_5_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_5_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_6_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_6_altOrBasePred;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_7_useProvider;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerTableIdx;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerWayIdx;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerTakenCtr_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerUsefulCtr_value;
    logic io_toFtq_meta_bits_resolveMeta_tage_entries_7_altOrBasePred;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_0;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_1;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_2;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_3;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_4;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_5;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_6;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_7;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_0;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_1;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_2;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_3;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_4;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_5;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_6;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_7;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_0;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_1;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_2;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_3;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_4;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_5;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_6;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_7;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_8;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_9;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_10;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_11;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_12;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_13;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_14;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_15;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_16;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_17;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_18;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_19;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_20;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_21;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_22;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_23;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_24;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_25;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_26;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_27;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_28;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_29;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_30;
    logic [5:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_31;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_0;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_1;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_2;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_3;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_4;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_5;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_6;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_valid;
    logic [15:0] io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_ghr;
    logic [7:0] io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_bw;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_scPred_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePred_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_useScPred_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_7;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_0;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_1;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_2;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_3;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_4;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_5;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_6;
    logic io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_7;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predPathIdx_0;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predPathIdx_1;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predGlobalIdx_0;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predGlobalIdx_1;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predBWIdx_0;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predBWIdx_1;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_sc_debug_predBiasIdx;
    logic io_toFtq_meta_bits_resolveMeta_ittage_provider_valid;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_ittage_provider_bits;
    logic io_toFtq_meta_bits_resolveMeta_ittage_altProvider_valid;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_ittage_altProvider_bits;
    logic io_toFtq_meta_bits_resolveMeta_ittage_altDiffers;
    logic io_toFtq_meta_bits_resolveMeta_ittage_providerUsefulCnt_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_ittage_providerCnt_value;
    logic [1:0] io_toFtq_meta_bits_resolveMeta_ittage_altProviderCnt_value;
    logic io_toFtq_meta_bits_resolveMeta_ittage_allocate_valid;
    logic [2:0] io_toFtq_meta_bits_resolveMeta_ittage_allocate_bits;
    logic [48:0] io_toFtq_meta_bits_resolveMeta_ittage_providerTarget_addr;
    logic [48:0] io_toFtq_meta_bits_resolveMeta_ittage_altProviderTarget_addr;
    logic [9:0] io_toFtq_meta_bits_resolveMeta_phr_phrPtr_value;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_phrLowBits;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_31_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_30_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_29_foldedHist;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_28_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_27_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_26_foldedHist;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_25_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_24_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_23_foldedHist;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_22_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_21_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_20_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_19_foldedHist;
    logic [7:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_18_foldedHist;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_17_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_16_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_15_foldedHist;
    logic [12:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_14_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_13_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_12_foldedHist;
    logic [11:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_11_foldedHist;
    logic [10:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_10_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_9_foldedHist;
    logic [7:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_8_foldedHist;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_7_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_6_foldedHist;
    logic [7:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_5_foldedHist;
    logic [8:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_4_foldedHist;
    logic [7:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_3_foldedHist;
    logic [7:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_2_foldedHist;
    logic [6:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_1_foldedHist;
    logic [3:0] io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_0_foldedHist;
    logic [3:0] io_toFtq_meta_bits_commitMeta_ras_ssp;
    logic io_toFtq_meta_bits_commitMeta_ras_tosw_flag;
    logic [4:0] io_toFtq_meta_bits_commitMeta_ras_tosw_value;
    logic io_toFtq_s3FtqPtr_flag;
    logic [5:0] io_toFtq_s3FtqPtr_value;
    logic [4:0] io_toFtq_perfMeta_s1Prediction_cfiPosition;
    logic [48:0] io_toFtq_perfMeta_s1Prediction_target_addr;
    logic [1:0] io_toFtq_perfMeta_s1Prediction_attribute_branchType;
    logic [1:0] io_toFtq_perfMeta_s1Prediction_attribute_rasAction;
    logic io_toFtq_perfMeta_s1Prediction_taken;
    logic [4:0] io_toFtq_perfMeta_s3Prediction_cfiPosition;
    logic [48:0] io_toFtq_perfMeta_s3Prediction_target_addr;
    logic [1:0] io_toFtq_perfMeta_s3Prediction_attribute_branchType;
    logic [1:0] io_toFtq_perfMeta_s3Prediction_attribute_rasAction;
    logic io_toFtq_perfMeta_s3Prediction_taken;
    logic io_toFtq_perfMeta_mbtbMeta_entries_0_0_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_0_0_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_0_1_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_0_1_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_0_2_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_0_2_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_0_3_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_0_3_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_1_0_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_1_0_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_1_1_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_1_1_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_1_2_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_1_2_position;
    logic io_toFtq_perfMeta_mbtbMeta_entries_1_3_rawHit;
    logic [4:0] io_toFtq_perfMeta_mbtbMeta_entries_1_3_position;
    logic [2:0] io_toFtq_perfMeta_bpSource_s1Source;
    logic [2:0] io_toFtq_perfMeta_bpSource_s3Source;
    logic io_toFtq_perfMeta_bpSource_s3Override;
    logic boreChildrenBd_bore_ack;
    logic [111:0] boreChildrenBd_bore_outdata;
    logic boreChildrenBd_bore_1_ack;
    logic [37:0] boreChildrenBd_bore_1_outdata;
    logic boreChildrenBd_bore_2_ack;
    logic [75:0] boreChildrenBd_bore_2_outdata;
    logic boreChildrenBd_bore_3_ack;
    logic [75:0] boreChildrenBd_bore_3_outdata;
    logic boreChildrenBd_bore_4_ack;
    logic [75:0] boreChildrenBd_bore_4_outdata;
    logic [47:0] boreChildrenBd_bore_5_rdata;
    logic [47:0] boreChildrenBd_bore_6_rdata;
    logic [47:0] boreChildrenBd_bore_7_rdata;
    logic [47:0] boreChildrenBd_bore_8_rdata;
    logic [47:0] boreChildrenBd_bore_9_rdata;
    logic [47:0] boreChildrenBd_bore_10_rdata;
    logic [47:0] boreChildrenBd_bore_11_rdata;
    logic [47:0] boreChildrenBd_bore_12_rdata;
    logic [47:0] boreChildrenBd_bore_13_rdata;
    logic [47:0] boreChildrenBd_bore_14_rdata;
    logic [47:0] boreChildrenBd_bore_15_rdata;
    logic [47:0] boreChildrenBd_bore_16_rdata;
    logic [191:0] boreChildrenBd_bore_17_rdata;
    logic [191:0] boreChildrenBd_bore_18_rdata;

    Bpu dut (
        .clock(clock),
        .reset(reset),
        .io_ctrl_ubtbEnable(io_ctrl_ubtbEnable),
        .io_ctrl_abtbEnable(io_ctrl_abtbEnable),
        .io_ctrl_mbtbEnable(io_ctrl_mbtbEnable),
        .io_ctrl_tageEnable(io_ctrl_tageEnable),
        .io_ctrl_scEnable(io_ctrl_scEnable),
        .io_ctrl_ittageEnable(io_ctrl_ittageEnable),
        .io_resetVector_addr(io_resetVector_addr),
        .io_fromFtq_redirect_valid(io_fromFtq_redirect_valid),
        .io_fromFtq_redirect_bits_cfiPc_addr(io_fromFtq_redirect_bits_cfiPc_addr),
        .io_fromFtq_redirect_bits_target_addr(io_fromFtq_redirect_bits_target_addr),
        .io_fromFtq_redirect_bits_taken(io_fromFtq_redirect_bits_taken),
        .io_fromFtq_redirect_bits_attribute_branchType(io_fromFtq_redirect_bits_attribute_branchType),
        .io_fromFtq_redirect_bits_attribute_rasAction(io_fromFtq_redirect_bits_attribute_rasAction),
        .io_fromFtq_redirect_bits_meta_phr_phrPtr_flag(io_fromFtq_redirect_bits_meta_phr_phrPtr_flag),
        .io_fromFtq_redirect_bits_meta_phr_phrPtr_value(io_fromFtq_redirect_bits_meta_phr_phrPtr_value),
        .io_fromFtq_redirect_bits_meta_phr_phrLowBits(io_fromFtq_redirect_bits_meta_phr_phrLowBits),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_ghr(io_fromFtq_redirect_bits_meta_commonHRMeta_ghr),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_bw(io_fromFtq_redirect_bits_meta_commonHRMeta_bw),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_0(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_0),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_1(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_1),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_2(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_2),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_3(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_3),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_4(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_4),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_5(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_5),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_6(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_6),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_7(io_fromFtq_redirect_bits_meta_commonHRMeta_hitMask_7),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_0_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_0_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_1_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_1_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_2_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_2_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_3_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_3_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_4_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_4_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_5_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_5_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_6_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_6_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_7_branchType(io_fromFtq_redirect_bits_meta_commonHRMeta_attribute_7_branchType),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_0(io_fromFtq_redirect_bits_meta_commonHRMeta_position_0),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_1(io_fromFtq_redirect_bits_meta_commonHRMeta_position_1),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_2(io_fromFtq_redirect_bits_meta_commonHRMeta_position_2),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_3(io_fromFtq_redirect_bits_meta_commonHRMeta_position_3),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_4(io_fromFtq_redirect_bits_meta_commonHRMeta_position_4),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_5(io_fromFtq_redirect_bits_meta_commonHRMeta_position_5),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_6(io_fromFtq_redirect_bits_meta_commonHRMeta_position_6),
        .io_fromFtq_redirect_bits_meta_commonHRMeta_position_7(io_fromFtq_redirect_bits_meta_commonHRMeta_position_7),
        .io_fromFtq_redirect_bits_meta_ras_ssp(io_fromFtq_redirect_bits_meta_ras_ssp),
        .io_fromFtq_redirect_bits_meta_ras_sctr(io_fromFtq_redirect_bits_meta_ras_sctr),
        .io_fromFtq_redirect_bits_meta_ras_tosw_flag(io_fromFtq_redirect_bits_meta_ras_tosw_flag),
        .io_fromFtq_redirect_bits_meta_ras_tosw_value(io_fromFtq_redirect_bits_meta_ras_tosw_value),
        .io_fromFtq_redirect_bits_meta_ras_tosr_flag(io_fromFtq_redirect_bits_meta_ras_tosr_flag),
        .io_fromFtq_redirect_bits_meta_ras_tosr_value(io_fromFtq_redirect_bits_meta_ras_tosr_value),
        .io_fromFtq_redirect_bits_meta_ras_nos_flag(io_fromFtq_redirect_bits_meta_ras_nos_flag),
        .io_fromFtq_redirect_bits_meta_ras_nos_value(io_fromFtq_redirect_bits_meta_ras_nos_value),
        .io_fromFtq_train_ready(io_fromFtq_train_ready),
        .io_fromFtq_train_valid(io_fromFtq_train_valid),
        .io_fromFtq_train_bits_startPc_addr(io_fromFtq_train_bits_startPc_addr),
        .io_fromFtq_train_bits_branches_0_valid(io_fromFtq_train_bits_branches_0_valid),
        .io_fromFtq_train_bits_branches_0_bits_target_addr(io_fromFtq_train_bits_branches_0_bits_target_addr),
        .io_fromFtq_train_bits_branches_0_bits_taken(io_fromFtq_train_bits_branches_0_bits_taken),
        .io_fromFtq_train_bits_branches_0_bits_cfiPosition(io_fromFtq_train_bits_branches_0_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_0_bits_attribute_branchType(io_fromFtq_train_bits_branches_0_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_0_bits_attribute_rasAction(io_fromFtq_train_bits_branches_0_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_0_bits_mispredict(io_fromFtq_train_bits_branches_0_bits_mispredict),
        .io_fromFtq_train_bits_branches_1_valid(io_fromFtq_train_bits_branches_1_valid),
        .io_fromFtq_train_bits_branches_1_bits_target_addr(io_fromFtq_train_bits_branches_1_bits_target_addr),
        .io_fromFtq_train_bits_branches_1_bits_taken(io_fromFtq_train_bits_branches_1_bits_taken),
        .io_fromFtq_train_bits_branches_1_bits_cfiPosition(io_fromFtq_train_bits_branches_1_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_1_bits_attribute_branchType(io_fromFtq_train_bits_branches_1_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_1_bits_attribute_rasAction(io_fromFtq_train_bits_branches_1_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_1_bits_mispredict(io_fromFtq_train_bits_branches_1_bits_mispredict),
        .io_fromFtq_train_bits_branches_2_valid(io_fromFtq_train_bits_branches_2_valid),
        .io_fromFtq_train_bits_branches_2_bits_target_addr(io_fromFtq_train_bits_branches_2_bits_target_addr),
        .io_fromFtq_train_bits_branches_2_bits_taken(io_fromFtq_train_bits_branches_2_bits_taken),
        .io_fromFtq_train_bits_branches_2_bits_cfiPosition(io_fromFtq_train_bits_branches_2_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_2_bits_attribute_branchType(io_fromFtq_train_bits_branches_2_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_2_bits_attribute_rasAction(io_fromFtq_train_bits_branches_2_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_2_bits_mispredict(io_fromFtq_train_bits_branches_2_bits_mispredict),
        .io_fromFtq_train_bits_branches_3_valid(io_fromFtq_train_bits_branches_3_valid),
        .io_fromFtq_train_bits_branches_3_bits_target_addr(io_fromFtq_train_bits_branches_3_bits_target_addr),
        .io_fromFtq_train_bits_branches_3_bits_taken(io_fromFtq_train_bits_branches_3_bits_taken),
        .io_fromFtq_train_bits_branches_3_bits_cfiPosition(io_fromFtq_train_bits_branches_3_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_3_bits_attribute_branchType(io_fromFtq_train_bits_branches_3_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_3_bits_attribute_rasAction(io_fromFtq_train_bits_branches_3_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_3_bits_mispredict(io_fromFtq_train_bits_branches_3_bits_mispredict),
        .io_fromFtq_train_bits_branches_4_valid(io_fromFtq_train_bits_branches_4_valid),
        .io_fromFtq_train_bits_branches_4_bits_target_addr(io_fromFtq_train_bits_branches_4_bits_target_addr),
        .io_fromFtq_train_bits_branches_4_bits_taken(io_fromFtq_train_bits_branches_4_bits_taken),
        .io_fromFtq_train_bits_branches_4_bits_cfiPosition(io_fromFtq_train_bits_branches_4_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_4_bits_attribute_branchType(io_fromFtq_train_bits_branches_4_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_4_bits_attribute_rasAction(io_fromFtq_train_bits_branches_4_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_4_bits_mispredict(io_fromFtq_train_bits_branches_4_bits_mispredict),
        .io_fromFtq_train_bits_branches_5_valid(io_fromFtq_train_bits_branches_5_valid),
        .io_fromFtq_train_bits_branches_5_bits_target_addr(io_fromFtq_train_bits_branches_5_bits_target_addr),
        .io_fromFtq_train_bits_branches_5_bits_taken(io_fromFtq_train_bits_branches_5_bits_taken),
        .io_fromFtq_train_bits_branches_5_bits_cfiPosition(io_fromFtq_train_bits_branches_5_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_5_bits_attribute_branchType(io_fromFtq_train_bits_branches_5_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_5_bits_attribute_rasAction(io_fromFtq_train_bits_branches_5_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_5_bits_mispredict(io_fromFtq_train_bits_branches_5_bits_mispredict),
        .io_fromFtq_train_bits_branches_6_valid(io_fromFtq_train_bits_branches_6_valid),
        .io_fromFtq_train_bits_branches_6_bits_target_addr(io_fromFtq_train_bits_branches_6_bits_target_addr),
        .io_fromFtq_train_bits_branches_6_bits_taken(io_fromFtq_train_bits_branches_6_bits_taken),
        .io_fromFtq_train_bits_branches_6_bits_cfiPosition(io_fromFtq_train_bits_branches_6_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_6_bits_attribute_branchType(io_fromFtq_train_bits_branches_6_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_6_bits_attribute_rasAction(io_fromFtq_train_bits_branches_6_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_6_bits_mispredict(io_fromFtq_train_bits_branches_6_bits_mispredict),
        .io_fromFtq_train_bits_branches_7_valid(io_fromFtq_train_bits_branches_7_valid),
        .io_fromFtq_train_bits_branches_7_bits_target_addr(io_fromFtq_train_bits_branches_7_bits_target_addr),
        .io_fromFtq_train_bits_branches_7_bits_taken(io_fromFtq_train_bits_branches_7_bits_taken),
        .io_fromFtq_train_bits_branches_7_bits_cfiPosition(io_fromFtq_train_bits_branches_7_bits_cfiPosition),
        .io_fromFtq_train_bits_branches_7_bits_attribute_branchType(io_fromFtq_train_bits_branches_7_bits_attribute_branchType),
        .io_fromFtq_train_bits_branches_7_bits_attribute_rasAction(io_fromFtq_train_bits_branches_7_bits_attribute_rasAction),
        .io_fromFtq_train_bits_branches_7_bits_mispredict(io_fromFtq_train_bits_branches_7_bits_mispredict),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_0_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_0_0_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_0_position(io_fromFtq_train_bits_meta_mbtb_entries_0_0_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_0_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_0_0_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_0_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_0_0_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_0_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_0_0_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_1_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_0_1_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_1_position(io_fromFtq_train_bits_meta_mbtb_entries_0_1_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_1_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_0_1_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_1_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_0_1_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_1_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_0_1_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_2_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_0_2_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_2_position(io_fromFtq_train_bits_meta_mbtb_entries_0_2_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_2_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_0_2_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_2_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_0_2_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_2_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_0_2_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_3_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_0_3_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_3_position(io_fromFtq_train_bits_meta_mbtb_entries_0_3_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_3_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_0_3_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_3_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_0_3_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_0_3_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_0_3_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_0_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_1_0_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_0_position(io_fromFtq_train_bits_meta_mbtb_entries_1_0_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_0_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_1_0_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_0_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_1_0_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_0_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_1_0_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_1_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_1_1_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_1_position(io_fromFtq_train_bits_meta_mbtb_entries_1_1_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_1_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_1_1_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_1_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_1_1_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_1_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_1_1_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_2_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_1_2_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_2_position(io_fromFtq_train_bits_meta_mbtb_entries_1_2_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_2_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_1_2_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_2_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_1_2_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_2_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_1_2_counter_value),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_3_rawHit(io_fromFtq_train_bits_meta_mbtb_entries_1_3_rawHit),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_3_position(io_fromFtq_train_bits_meta_mbtb_entries_1_3_position),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_3_attribute_branchType(io_fromFtq_train_bits_meta_mbtb_entries_1_3_attribute_branchType),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_3_attribute_rasAction(io_fromFtq_train_bits_meta_mbtb_entries_1_3_attribute_rasAction),
        .io_fromFtq_train_bits_meta_mbtb_entries_1_3_counter_value(io_fromFtq_train_bits_meta_mbtb_entries_1_3_counter_value),
        .io_fromFtq_train_bits_meta_tage_entries_0_useProvider(io_fromFtq_train_bits_meta_tage_entries_0_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_0_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_0_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_0_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_0_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_0_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_0_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_0_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_0_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_0_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_0_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_1_useProvider(io_fromFtq_train_bits_meta_tage_entries_1_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_1_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_1_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_1_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_1_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_1_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_1_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_1_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_1_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_1_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_1_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_2_useProvider(io_fromFtq_train_bits_meta_tage_entries_2_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_2_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_2_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_2_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_2_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_2_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_2_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_2_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_2_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_2_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_2_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_3_useProvider(io_fromFtq_train_bits_meta_tage_entries_3_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_3_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_3_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_3_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_3_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_3_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_3_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_3_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_3_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_3_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_3_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_4_useProvider(io_fromFtq_train_bits_meta_tage_entries_4_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_4_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_4_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_4_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_4_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_4_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_4_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_4_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_4_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_4_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_4_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_5_useProvider(io_fromFtq_train_bits_meta_tage_entries_5_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_5_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_5_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_5_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_5_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_5_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_5_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_5_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_5_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_5_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_5_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_6_useProvider(io_fromFtq_train_bits_meta_tage_entries_6_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_6_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_6_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_6_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_6_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_6_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_6_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_6_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_6_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_6_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_6_altOrBasePred),
        .io_fromFtq_train_bits_meta_tage_entries_7_useProvider(io_fromFtq_train_bits_meta_tage_entries_7_useProvider),
        .io_fromFtq_train_bits_meta_tage_entries_7_providerTableIdx(io_fromFtq_train_bits_meta_tage_entries_7_providerTableIdx),
        .io_fromFtq_train_bits_meta_tage_entries_7_providerWayIdx(io_fromFtq_train_bits_meta_tage_entries_7_providerWayIdx),
        .io_fromFtq_train_bits_meta_tage_entries_7_providerTakenCtr_value(io_fromFtq_train_bits_meta_tage_entries_7_providerTakenCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_7_providerUsefulCtr_value(io_fromFtq_train_bits_meta_tage_entries_7_providerUsefulCtr_value),
        .io_fromFtq_train_bits_meta_tage_entries_7_altOrBasePred(io_fromFtq_train_bits_meta_tage_entries_7_altOrBasePred),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_0(io_fromFtq_train_bits_meta_sc_scPathResp_0_0),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_1(io_fromFtq_train_bits_meta_sc_scPathResp_0_1),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_2(io_fromFtq_train_bits_meta_sc_scPathResp_0_2),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_3(io_fromFtq_train_bits_meta_sc_scPathResp_0_3),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_4(io_fromFtq_train_bits_meta_sc_scPathResp_0_4),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_5(io_fromFtq_train_bits_meta_sc_scPathResp_0_5),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_6(io_fromFtq_train_bits_meta_sc_scPathResp_0_6),
        .io_fromFtq_train_bits_meta_sc_scPathResp_0_7(io_fromFtq_train_bits_meta_sc_scPathResp_0_7),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_0(io_fromFtq_train_bits_meta_sc_scPathResp_1_0),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_1(io_fromFtq_train_bits_meta_sc_scPathResp_1_1),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_2(io_fromFtq_train_bits_meta_sc_scPathResp_1_2),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_3(io_fromFtq_train_bits_meta_sc_scPathResp_1_3),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_4(io_fromFtq_train_bits_meta_sc_scPathResp_1_4),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_5(io_fromFtq_train_bits_meta_sc_scPathResp_1_5),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_6(io_fromFtq_train_bits_meta_sc_scPathResp_1_6),
        .io_fromFtq_train_bits_meta_sc_scPathResp_1_7(io_fromFtq_train_bits_meta_sc_scPathResp_1_7),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_0(io_fromFtq_train_bits_meta_sc_scBiasResp_0),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_1(io_fromFtq_train_bits_meta_sc_scBiasResp_1),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_2(io_fromFtq_train_bits_meta_sc_scBiasResp_2),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_3(io_fromFtq_train_bits_meta_sc_scBiasResp_3),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_4(io_fromFtq_train_bits_meta_sc_scBiasResp_4),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_5(io_fromFtq_train_bits_meta_sc_scBiasResp_5),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_6(io_fromFtq_train_bits_meta_sc_scBiasResp_6),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_7(io_fromFtq_train_bits_meta_sc_scBiasResp_7),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_8(io_fromFtq_train_bits_meta_sc_scBiasResp_8),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_9(io_fromFtq_train_bits_meta_sc_scBiasResp_9),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_10(io_fromFtq_train_bits_meta_sc_scBiasResp_10),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_11(io_fromFtq_train_bits_meta_sc_scBiasResp_11),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_12(io_fromFtq_train_bits_meta_sc_scBiasResp_12),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_13(io_fromFtq_train_bits_meta_sc_scBiasResp_13),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_14(io_fromFtq_train_bits_meta_sc_scBiasResp_14),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_15(io_fromFtq_train_bits_meta_sc_scBiasResp_15),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_16(io_fromFtq_train_bits_meta_sc_scBiasResp_16),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_17(io_fromFtq_train_bits_meta_sc_scBiasResp_17),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_18(io_fromFtq_train_bits_meta_sc_scBiasResp_18),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_19(io_fromFtq_train_bits_meta_sc_scBiasResp_19),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_20(io_fromFtq_train_bits_meta_sc_scBiasResp_20),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_21(io_fromFtq_train_bits_meta_sc_scBiasResp_21),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_22(io_fromFtq_train_bits_meta_sc_scBiasResp_22),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_23(io_fromFtq_train_bits_meta_sc_scBiasResp_23),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_24(io_fromFtq_train_bits_meta_sc_scBiasResp_24),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_25(io_fromFtq_train_bits_meta_sc_scBiasResp_25),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_26(io_fromFtq_train_bits_meta_sc_scBiasResp_26),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_27(io_fromFtq_train_bits_meta_sc_scBiasResp_27),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_28(io_fromFtq_train_bits_meta_sc_scBiasResp_28),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_29(io_fromFtq_train_bits_meta_sc_scBiasResp_29),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_30(io_fromFtq_train_bits_meta_sc_scBiasResp_30),
        .io_fromFtq_train_bits_meta_sc_scBiasResp_31(io_fromFtq_train_bits_meta_sc_scBiasResp_31),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_0(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_0),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_1(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_1),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_2(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_2),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_3(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_3),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_4(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_4),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_5(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_5),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_6(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_6),
        .io_fromFtq_train_bits_meta_sc_scBiasLowerBits_7(io_fromFtq_train_bits_meta_sc_scBiasLowerBits_7),
        .io_fromFtq_train_bits_meta_sc_scCommonHR_valid(io_fromFtq_train_bits_meta_sc_scCommonHR_valid),
        .io_fromFtq_train_bits_meta_sc_scCommonHR_ghr(io_fromFtq_train_bits_meta_sc_scCommonHR_ghr),
        .io_fromFtq_train_bits_meta_sc_scCommonHR_bw(io_fromFtq_train_bits_meta_sc_scCommonHR_bw),
        .io_fromFtq_train_bits_meta_sc_scPred_0(io_fromFtq_train_bits_meta_sc_scPred_0),
        .io_fromFtq_train_bits_meta_sc_scPred_1(io_fromFtq_train_bits_meta_sc_scPred_1),
        .io_fromFtq_train_bits_meta_sc_scPred_2(io_fromFtq_train_bits_meta_sc_scPred_2),
        .io_fromFtq_train_bits_meta_sc_scPred_3(io_fromFtq_train_bits_meta_sc_scPred_3),
        .io_fromFtq_train_bits_meta_sc_scPred_4(io_fromFtq_train_bits_meta_sc_scPred_4),
        .io_fromFtq_train_bits_meta_sc_scPred_5(io_fromFtq_train_bits_meta_sc_scPred_5),
        .io_fromFtq_train_bits_meta_sc_scPred_6(io_fromFtq_train_bits_meta_sc_scPred_6),
        .io_fromFtq_train_bits_meta_sc_scPred_7(io_fromFtq_train_bits_meta_sc_scPred_7),
        .io_fromFtq_train_bits_meta_sc_tagePred_0(io_fromFtq_train_bits_meta_sc_tagePred_0),
        .io_fromFtq_train_bits_meta_sc_tagePred_1(io_fromFtq_train_bits_meta_sc_tagePred_1),
        .io_fromFtq_train_bits_meta_sc_tagePred_2(io_fromFtq_train_bits_meta_sc_tagePred_2),
        .io_fromFtq_train_bits_meta_sc_tagePred_3(io_fromFtq_train_bits_meta_sc_tagePred_3),
        .io_fromFtq_train_bits_meta_sc_tagePred_4(io_fromFtq_train_bits_meta_sc_tagePred_4),
        .io_fromFtq_train_bits_meta_sc_tagePred_5(io_fromFtq_train_bits_meta_sc_tagePred_5),
        .io_fromFtq_train_bits_meta_sc_tagePred_6(io_fromFtq_train_bits_meta_sc_tagePred_6),
        .io_fromFtq_train_bits_meta_sc_tagePred_7(io_fromFtq_train_bits_meta_sc_tagePred_7),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_0(io_fromFtq_train_bits_meta_sc_tagePredValid_0),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_1(io_fromFtq_train_bits_meta_sc_tagePredValid_1),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_2(io_fromFtq_train_bits_meta_sc_tagePredValid_2),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_3(io_fromFtq_train_bits_meta_sc_tagePredValid_3),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_4(io_fromFtq_train_bits_meta_sc_tagePredValid_4),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_5(io_fromFtq_train_bits_meta_sc_tagePredValid_5),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_6(io_fromFtq_train_bits_meta_sc_tagePredValid_6),
        .io_fromFtq_train_bits_meta_sc_tagePredValid_7(io_fromFtq_train_bits_meta_sc_tagePredValid_7),
        .io_fromFtq_train_bits_meta_sc_useScPred_0(io_fromFtq_train_bits_meta_sc_useScPred_0),
        .io_fromFtq_train_bits_meta_sc_useScPred_1(io_fromFtq_train_bits_meta_sc_useScPred_1),
        .io_fromFtq_train_bits_meta_sc_useScPred_2(io_fromFtq_train_bits_meta_sc_useScPred_2),
        .io_fromFtq_train_bits_meta_sc_useScPred_3(io_fromFtq_train_bits_meta_sc_useScPred_3),
        .io_fromFtq_train_bits_meta_sc_useScPred_4(io_fromFtq_train_bits_meta_sc_useScPred_4),
        .io_fromFtq_train_bits_meta_sc_useScPred_5(io_fromFtq_train_bits_meta_sc_useScPred_5),
        .io_fromFtq_train_bits_meta_sc_useScPred_6(io_fromFtq_train_bits_meta_sc_useScPred_6),
        .io_fromFtq_train_bits_meta_sc_useScPred_7(io_fromFtq_train_bits_meta_sc_useScPred_7),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_0(io_fromFtq_train_bits_meta_sc_sumAboveThres_0),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_1(io_fromFtq_train_bits_meta_sc_sumAboveThres_1),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_2(io_fromFtq_train_bits_meta_sc_sumAboveThres_2),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_3(io_fromFtq_train_bits_meta_sc_sumAboveThres_3),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_4(io_fromFtq_train_bits_meta_sc_sumAboveThres_4),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_5(io_fromFtq_train_bits_meta_sc_sumAboveThres_5),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_6(io_fromFtq_train_bits_meta_sc_sumAboveThres_6),
        .io_fromFtq_train_bits_meta_sc_sumAboveThres_7(io_fromFtq_train_bits_meta_sc_sumAboveThres_7),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_0(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_0),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_1(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_1),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_2(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_2),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_3(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_3),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_4(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_4),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_5(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_5),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_6(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_6),
        .io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_7(io_fromFtq_train_bits_meta_sc_debug_scPathTakenVec_7),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_0(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_0),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_1(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_1),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_2(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_2),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_3(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_3),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_4(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_4),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_5(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_5),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_6(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_6),
        .io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_7(io_fromFtq_train_bits_meta_sc_debug_scBiasTakenVec_7),
        .io_fromFtq_train_bits_meta_sc_debug_predPathIdx_0(io_fromFtq_train_bits_meta_sc_debug_predPathIdx_0),
        .io_fromFtq_train_bits_meta_sc_debug_predPathIdx_1(io_fromFtq_train_bits_meta_sc_debug_predPathIdx_1),
        .io_fromFtq_train_bits_meta_sc_debug_predGlobalIdx_0(io_fromFtq_train_bits_meta_sc_debug_predGlobalIdx_0),
        .io_fromFtq_train_bits_meta_sc_debug_predGlobalIdx_1(io_fromFtq_train_bits_meta_sc_debug_predGlobalIdx_1),
        .io_fromFtq_train_bits_meta_sc_debug_predBWIdx_0(io_fromFtq_train_bits_meta_sc_debug_predBWIdx_0),
        .io_fromFtq_train_bits_meta_sc_debug_predBWIdx_1(io_fromFtq_train_bits_meta_sc_debug_predBWIdx_1),
        .io_fromFtq_train_bits_meta_sc_debug_predBiasIdx(io_fromFtq_train_bits_meta_sc_debug_predBiasIdx),
        .io_fromFtq_train_bits_meta_ittage_provider_valid(io_fromFtq_train_bits_meta_ittage_provider_valid),
        .io_fromFtq_train_bits_meta_ittage_provider_bits(io_fromFtq_train_bits_meta_ittage_provider_bits),
        .io_fromFtq_train_bits_meta_ittage_altProvider_valid(io_fromFtq_train_bits_meta_ittage_altProvider_valid),
        .io_fromFtq_train_bits_meta_ittage_altProvider_bits(io_fromFtq_train_bits_meta_ittage_altProvider_bits),
        .io_fromFtq_train_bits_meta_ittage_altDiffers(io_fromFtq_train_bits_meta_ittage_altDiffers),
        .io_fromFtq_train_bits_meta_ittage_providerUsefulCnt_value(io_fromFtq_train_bits_meta_ittage_providerUsefulCnt_value),
        .io_fromFtq_train_bits_meta_ittage_providerCnt_value(io_fromFtq_train_bits_meta_ittage_providerCnt_value),
        .io_fromFtq_train_bits_meta_ittage_altProviderCnt_value(io_fromFtq_train_bits_meta_ittage_altProviderCnt_value),
        .io_fromFtq_train_bits_meta_ittage_allocate_valid(io_fromFtq_train_bits_meta_ittage_allocate_valid),
        .io_fromFtq_train_bits_meta_ittage_allocate_bits(io_fromFtq_train_bits_meta_ittage_allocate_bits),
        .io_fromFtq_train_bits_meta_ittage_providerTarget_addr(io_fromFtq_train_bits_meta_ittage_providerTarget_addr),
        .io_fromFtq_train_bits_meta_ittage_altProviderTarget_addr(io_fromFtq_train_bits_meta_ittage_altProviderTarget_addr),
        .io_fromFtq_train_bits_meta_phr_phrPtr_value(io_fromFtq_train_bits_meta_phr_phrPtr_value),
        .io_fromFtq_train_bits_meta_phr_phrLowBits(io_fromFtq_train_bits_meta_phr_phrLowBits),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_31_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_31_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_30_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_30_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_29_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_29_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_28_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_28_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_27_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_27_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_26_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_26_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_25_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_25_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_24_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_24_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_23_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_23_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_22_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_22_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_21_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_21_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_20_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_20_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_19_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_19_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_18_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_18_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_17_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_17_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_16_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_16_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_15_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_15_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_14_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_14_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_13_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_13_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_12_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_12_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_11_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_11_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_10_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_10_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_9_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_9_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_8_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_8_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_7_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_7_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_6_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_6_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_5_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_5_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_4_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_4_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_3_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_3_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_2_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_2_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_1_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_1_foldedHist),
        .io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_0_foldedHist(io_fromFtq_train_bits_meta_phr_predFoldedHist_hist_0_foldedHist),
        .io_fromFtq_commit_valid(io_fromFtq_commit_valid),
        .io_fromFtq_commit_bits_meta_ras_ssp(io_fromFtq_commit_bits_meta_ras_ssp),
        .io_fromFtq_commit_bits_meta_ras_tosw_flag(io_fromFtq_commit_bits_meta_ras_tosw_flag),
        .io_fromFtq_commit_bits_meta_ras_tosw_value(io_fromFtq_commit_bits_meta_ras_tosw_value),
        .io_fromFtq_commit_bits_attribute_rasAction(io_fromFtq_commit_bits_attribute_rasAction),
        .io_fromFtq_bpuPtr_flag(io_fromFtq_bpuPtr_flag),
        .io_fromFtq_bpuPtr_value(io_fromFtq_bpuPtr_value),
        .io_toFtq_prediction_ready(io_toFtq_prediction_ready),
        .io_toFtq_prediction_valid(io_toFtq_prediction_valid),
        .io_toFtq_prediction_bits_startPc_addr(io_toFtq_prediction_bits_startPc_addr),
        .io_toFtq_prediction_bits_target_addr(io_toFtq_prediction_bits_target_addr),
        .io_toFtq_prediction_bits_takenCfiOffset_valid(io_toFtq_prediction_bits_takenCfiOffset_valid),
        .io_toFtq_prediction_bits_takenCfiOffset_bits(io_toFtq_prediction_bits_takenCfiOffset_bits),
        .io_toFtq_prediction_bits_s3Override(io_toFtq_prediction_bits_s3Override),
        .io_toFtq_meta_valid(io_toFtq_meta_valid),
        .io_toFtq_meta_bits_redirectMeta_phr_phrPtr_flag(io_toFtq_meta_bits_redirectMeta_phr_phrPtr_flag),
        .io_toFtq_meta_bits_redirectMeta_phr_phrPtr_value(io_toFtq_meta_bits_redirectMeta_phr_phrPtr_value),
        .io_toFtq_meta_bits_redirectMeta_phr_phrLowBits(io_toFtq_meta_bits_redirectMeta_phr_phrLowBits),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_ghr(io_toFtq_meta_bits_redirectMeta_commonHRMeta_ghr),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_bw(io_toFtq_meta_bits_redirectMeta_commonHRMeta_bw),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_0(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_0),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_1(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_1),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_2(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_2),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_3(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_3),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_4(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_4),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_5(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_5),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_6(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_6),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_7(io_toFtq_meta_bits_redirectMeta_commonHRMeta_hitMask_7),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_0_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_0_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_1_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_1_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_2_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_2_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_3_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_3_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_4_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_4_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_5_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_5_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_6_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_6_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_7_branchType(io_toFtq_meta_bits_redirectMeta_commonHRMeta_attribute_7_branchType),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_0(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_0),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_1(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_1),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_2(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_2),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_3(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_3),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_4(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_4),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_5(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_5),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_6(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_6),
        .io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_7(io_toFtq_meta_bits_redirectMeta_commonHRMeta_position_7),
        .io_toFtq_meta_bits_redirectMeta_ras_ssp(io_toFtq_meta_bits_redirectMeta_ras_ssp),
        .io_toFtq_meta_bits_redirectMeta_ras_sctr(io_toFtq_meta_bits_redirectMeta_ras_sctr),
        .io_toFtq_meta_bits_redirectMeta_ras_tosw_flag(io_toFtq_meta_bits_redirectMeta_ras_tosw_flag),
        .io_toFtq_meta_bits_redirectMeta_ras_tosw_value(io_toFtq_meta_bits_redirectMeta_ras_tosw_value),
        .io_toFtq_meta_bits_redirectMeta_ras_tosr_flag(io_toFtq_meta_bits_redirectMeta_ras_tosr_flag),
        .io_toFtq_meta_bits_redirectMeta_ras_tosr_value(io_toFtq_meta_bits_redirectMeta_ras_tosr_value),
        .io_toFtq_meta_bits_redirectMeta_ras_nos_flag(io_toFtq_meta_bits_redirectMeta_ras_nos_flag),
        .io_toFtq_meta_bits_redirectMeta_ras_nos_value(io_toFtq_meta_bits_redirectMeta_ras_nos_value),
        .io_toFtq_meta_bits_redirectMeta_ras_topRetAddr_addr(io_toFtq_meta_bits_redirectMeta_ras_topRetAddr_addr),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_0_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_1_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_2_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_0_3_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_0_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_1_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_2_counter_value),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_rawHit(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_rawHit),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_position(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_position),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_attribute_branchType(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_attribute_branchType),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_attribute_rasAction(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_attribute_rasAction),
        .io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_counter_value(io_toFtq_meta_bits_resolveMeta_mbtb_entries_1_3_counter_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_0_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_0_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_0_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_0_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_0_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_1_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_1_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_1_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_1_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_1_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_2_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_2_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_2_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_2_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_2_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_3_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_3_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_3_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_3_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_3_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_4_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_4_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_4_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_4_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_4_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_5_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_5_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_5_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_5_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_5_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_6_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_6_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_6_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_6_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_6_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_7_useProvider(io_toFtq_meta_bits_resolveMeta_tage_entries_7_useProvider),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerTableIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerTableIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerWayIdx(io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerWayIdx),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerTakenCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerTakenCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerUsefulCtr_value(io_toFtq_meta_bits_resolveMeta_tage_entries_7_providerUsefulCtr_value),
        .io_toFtq_meta_bits_resolveMeta_tage_entries_7_altOrBasePred(io_toFtq_meta_bits_resolveMeta_tage_entries_7_altOrBasePred),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_0(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_0),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_1(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_1),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_2(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_2),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_3(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_3),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_4(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_4),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_5(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_5),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_6(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_6),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_7(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_0_7),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_0(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_0),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_1(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_1),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_2(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_2),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_3(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_3),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_4(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_4),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_5(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_5),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_6(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_6),
        .io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_7(io_toFtq_meta_bits_resolveMeta_sc_scPathResp_1_7),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_0(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_0),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_1(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_1),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_2(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_2),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_3(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_3),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_4(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_4),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_5(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_5),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_6(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_6),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_7(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_7),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_8(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_8),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_9(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_9),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_10(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_10),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_11(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_11),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_12(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_12),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_13(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_13),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_14(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_14),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_15(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_15),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_16(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_16),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_17(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_17),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_18(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_18),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_19(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_19),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_20(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_20),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_21(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_21),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_22(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_22),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_23(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_23),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_24(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_24),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_25(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_25),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_26(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_26),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_27(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_27),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_28(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_28),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_29(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_29),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_30(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_30),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_31(io_toFtq_meta_bits_resolveMeta_sc_scBiasResp_31),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_0(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_0),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_1(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_1),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_2(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_2),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_3(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_3),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_4(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_4),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_5(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_5),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_6(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_6),
        .io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_7(io_toFtq_meta_bits_resolveMeta_sc_scBiasLowerBits_7),
        .io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_valid(io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_valid),
        .io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_ghr(io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_ghr),
        .io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_bw(io_toFtq_meta_bits_resolveMeta_sc_scCommonHR_bw),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_0(io_toFtq_meta_bits_resolveMeta_sc_scPred_0),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_1(io_toFtq_meta_bits_resolveMeta_sc_scPred_1),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_2(io_toFtq_meta_bits_resolveMeta_sc_scPred_2),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_3(io_toFtq_meta_bits_resolveMeta_sc_scPred_3),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_4(io_toFtq_meta_bits_resolveMeta_sc_scPred_4),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_5(io_toFtq_meta_bits_resolveMeta_sc_scPred_5),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_6(io_toFtq_meta_bits_resolveMeta_sc_scPred_6),
        .io_toFtq_meta_bits_resolveMeta_sc_scPred_7(io_toFtq_meta_bits_resolveMeta_sc_scPred_7),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_0(io_toFtq_meta_bits_resolveMeta_sc_tagePred_0),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_1(io_toFtq_meta_bits_resolveMeta_sc_tagePred_1),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_2(io_toFtq_meta_bits_resolveMeta_sc_tagePred_2),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_3(io_toFtq_meta_bits_resolveMeta_sc_tagePred_3),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_4(io_toFtq_meta_bits_resolveMeta_sc_tagePred_4),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_5(io_toFtq_meta_bits_resolveMeta_sc_tagePred_5),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_6(io_toFtq_meta_bits_resolveMeta_sc_tagePred_6),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePred_7(io_toFtq_meta_bits_resolveMeta_sc_tagePred_7),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_0(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_0),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_1(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_1),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_2(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_2),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_3(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_3),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_4(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_4),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_5(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_5),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_6(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_6),
        .io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_7(io_toFtq_meta_bits_resolveMeta_sc_tagePredValid_7),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_0(io_toFtq_meta_bits_resolveMeta_sc_useScPred_0),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_1(io_toFtq_meta_bits_resolveMeta_sc_useScPred_1),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_2(io_toFtq_meta_bits_resolveMeta_sc_useScPred_2),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_3(io_toFtq_meta_bits_resolveMeta_sc_useScPred_3),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_4(io_toFtq_meta_bits_resolveMeta_sc_useScPred_4),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_5(io_toFtq_meta_bits_resolveMeta_sc_useScPred_5),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_6(io_toFtq_meta_bits_resolveMeta_sc_useScPred_6),
        .io_toFtq_meta_bits_resolveMeta_sc_useScPred_7(io_toFtq_meta_bits_resolveMeta_sc_useScPred_7),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_0(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_0),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_1(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_1),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_2(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_2),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_3(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_3),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_4(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_4),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_5(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_5),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_6(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_6),
        .io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_7(io_toFtq_meta_bits_resolveMeta_sc_sumAboveThres_7),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_0(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_0),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_1(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_1),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_2(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_2),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_3(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_3),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_4(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_4),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_5(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_5),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_6(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_6),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_7(io_toFtq_meta_bits_resolveMeta_sc_debug_scPathTakenVec_7),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_0(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_0),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_1(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_1),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_2(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_2),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_3(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_3),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_4(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_4),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_5(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_5),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_6(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_6),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_7(io_toFtq_meta_bits_resolveMeta_sc_debug_scBiasTakenVec_7),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predPathIdx_0(io_toFtq_meta_bits_resolveMeta_sc_debug_predPathIdx_0),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predPathIdx_1(io_toFtq_meta_bits_resolveMeta_sc_debug_predPathIdx_1),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predGlobalIdx_0(io_toFtq_meta_bits_resolveMeta_sc_debug_predGlobalIdx_0),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predGlobalIdx_1(io_toFtq_meta_bits_resolveMeta_sc_debug_predGlobalIdx_1),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predBWIdx_0(io_toFtq_meta_bits_resolveMeta_sc_debug_predBWIdx_0),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predBWIdx_1(io_toFtq_meta_bits_resolveMeta_sc_debug_predBWIdx_1),
        .io_toFtq_meta_bits_resolveMeta_sc_debug_predBiasIdx(io_toFtq_meta_bits_resolveMeta_sc_debug_predBiasIdx),
        .io_toFtq_meta_bits_resolveMeta_ittage_provider_valid(io_toFtq_meta_bits_resolveMeta_ittage_provider_valid),
        .io_toFtq_meta_bits_resolveMeta_ittage_provider_bits(io_toFtq_meta_bits_resolveMeta_ittage_provider_bits),
        .io_toFtq_meta_bits_resolveMeta_ittage_altProvider_valid(io_toFtq_meta_bits_resolveMeta_ittage_altProvider_valid),
        .io_toFtq_meta_bits_resolveMeta_ittage_altProvider_bits(io_toFtq_meta_bits_resolveMeta_ittage_altProvider_bits),
        .io_toFtq_meta_bits_resolveMeta_ittage_altDiffers(io_toFtq_meta_bits_resolveMeta_ittage_altDiffers),
        .io_toFtq_meta_bits_resolveMeta_ittage_providerUsefulCnt_value(io_toFtq_meta_bits_resolveMeta_ittage_providerUsefulCnt_value),
        .io_toFtq_meta_bits_resolveMeta_ittage_providerCnt_value(io_toFtq_meta_bits_resolveMeta_ittage_providerCnt_value),
        .io_toFtq_meta_bits_resolveMeta_ittage_altProviderCnt_value(io_toFtq_meta_bits_resolveMeta_ittage_altProviderCnt_value),
        .io_toFtq_meta_bits_resolveMeta_ittage_allocate_valid(io_toFtq_meta_bits_resolveMeta_ittage_allocate_valid),
        .io_toFtq_meta_bits_resolveMeta_ittage_allocate_bits(io_toFtq_meta_bits_resolveMeta_ittage_allocate_bits),
        .io_toFtq_meta_bits_resolveMeta_ittage_providerTarget_addr(io_toFtq_meta_bits_resolveMeta_ittage_providerTarget_addr),
        .io_toFtq_meta_bits_resolveMeta_ittage_altProviderTarget_addr(io_toFtq_meta_bits_resolveMeta_ittage_altProviderTarget_addr),
        .io_toFtq_meta_bits_resolveMeta_phr_phrPtr_value(io_toFtq_meta_bits_resolveMeta_phr_phrPtr_value),
        .io_toFtq_meta_bits_resolveMeta_phr_phrLowBits(io_toFtq_meta_bits_resolveMeta_phr_phrLowBits),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_31_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_31_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_30_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_30_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_29_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_29_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_28_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_28_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_27_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_27_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_26_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_26_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_25_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_25_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_24_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_24_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_23_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_23_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_22_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_22_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_21_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_21_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_20_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_20_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_19_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_19_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_18_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_18_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_17_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_17_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_16_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_16_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_15_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_15_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_14_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_14_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_13_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_13_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_12_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_12_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_11_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_11_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_10_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_10_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_9_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_9_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_8_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_8_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_7_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_7_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_6_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_6_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_5_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_5_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_4_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_4_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_3_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_3_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_2_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_2_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_1_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_1_foldedHist),
        .io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_0_foldedHist(io_toFtq_meta_bits_resolveMeta_phr_predFoldedHist_hist_0_foldedHist),
        .io_toFtq_meta_bits_commitMeta_ras_ssp(io_toFtq_meta_bits_commitMeta_ras_ssp),
        .io_toFtq_meta_bits_commitMeta_ras_tosw_flag(io_toFtq_meta_bits_commitMeta_ras_tosw_flag),
        .io_toFtq_meta_bits_commitMeta_ras_tosw_value(io_toFtq_meta_bits_commitMeta_ras_tosw_value),
        .io_toFtq_s3FtqPtr_flag(io_toFtq_s3FtqPtr_flag),
        .io_toFtq_s3FtqPtr_value(io_toFtq_s3FtqPtr_value),
        .io_toFtq_perfMeta_s1Prediction_cfiPosition(io_toFtq_perfMeta_s1Prediction_cfiPosition),
        .io_toFtq_perfMeta_s1Prediction_target_addr(io_toFtq_perfMeta_s1Prediction_target_addr),
        .io_toFtq_perfMeta_s1Prediction_attribute_branchType(io_toFtq_perfMeta_s1Prediction_attribute_branchType),
        .io_toFtq_perfMeta_s1Prediction_attribute_rasAction(io_toFtq_perfMeta_s1Prediction_attribute_rasAction),
        .io_toFtq_perfMeta_s1Prediction_taken(io_toFtq_perfMeta_s1Prediction_taken),
        .io_toFtq_perfMeta_s3Prediction_cfiPosition(io_toFtq_perfMeta_s3Prediction_cfiPosition),
        .io_toFtq_perfMeta_s3Prediction_target_addr(io_toFtq_perfMeta_s3Prediction_target_addr),
        .io_toFtq_perfMeta_s3Prediction_attribute_branchType(io_toFtq_perfMeta_s3Prediction_attribute_branchType),
        .io_toFtq_perfMeta_s3Prediction_attribute_rasAction(io_toFtq_perfMeta_s3Prediction_attribute_rasAction),
        .io_toFtq_perfMeta_s3Prediction_taken(io_toFtq_perfMeta_s3Prediction_taken),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_0_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_0_0_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_0_position(io_toFtq_perfMeta_mbtbMeta_entries_0_0_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_1_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_0_1_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_1_position(io_toFtq_perfMeta_mbtbMeta_entries_0_1_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_2_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_0_2_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_2_position(io_toFtq_perfMeta_mbtbMeta_entries_0_2_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_3_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_0_3_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_0_3_position(io_toFtq_perfMeta_mbtbMeta_entries_0_3_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_0_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_1_0_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_0_position(io_toFtq_perfMeta_mbtbMeta_entries_1_0_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_1_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_1_1_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_1_position(io_toFtq_perfMeta_mbtbMeta_entries_1_1_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_2_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_1_2_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_2_position(io_toFtq_perfMeta_mbtbMeta_entries_1_2_position),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_3_rawHit(io_toFtq_perfMeta_mbtbMeta_entries_1_3_rawHit),
        .io_toFtq_perfMeta_mbtbMeta_entries_1_3_position(io_toFtq_perfMeta_mbtbMeta_entries_1_3_position),
        .io_toFtq_perfMeta_bpSource_s1Source(io_toFtq_perfMeta_bpSource_s1Source),
        .io_toFtq_perfMeta_bpSource_s3Source(io_toFtq_perfMeta_bpSource_s3Source),
        .io_toFtq_perfMeta_bpSource_s3Override(io_toFtq_perfMeta_bpSource_s3Override),
        .boreChildrenBd_bore_array(boreChildrenBd_bore_array),
        .boreChildrenBd_bore_all(boreChildrenBd_bore_all),
        .boreChildrenBd_bore_req(boreChildrenBd_bore_req),
        .boreChildrenBd_bore_ack(boreChildrenBd_bore_ack),
        .boreChildrenBd_bore_writeen(boreChildrenBd_bore_writeen),
        .boreChildrenBd_bore_be(boreChildrenBd_bore_be),
        .boreChildrenBd_bore_addr(boreChildrenBd_bore_addr),
        .boreChildrenBd_bore_indata(boreChildrenBd_bore_indata),
        .boreChildrenBd_bore_readen(boreChildrenBd_bore_readen),
        .boreChildrenBd_bore_addr_rd(boreChildrenBd_bore_addr_rd),
        .boreChildrenBd_bore_outdata(boreChildrenBd_bore_outdata),
        .boreChildrenBd_bore_1_array(boreChildrenBd_bore_1_array),
        .boreChildrenBd_bore_1_all(boreChildrenBd_bore_1_all),
        .boreChildrenBd_bore_1_req(boreChildrenBd_bore_1_req),
        .boreChildrenBd_bore_1_ack(boreChildrenBd_bore_1_ack),
        .boreChildrenBd_bore_1_writeen(boreChildrenBd_bore_1_writeen),
        .boreChildrenBd_bore_1_be(boreChildrenBd_bore_1_be),
        .boreChildrenBd_bore_1_addr(boreChildrenBd_bore_1_addr),
        .boreChildrenBd_bore_1_indata(boreChildrenBd_bore_1_indata),
        .boreChildrenBd_bore_1_readen(boreChildrenBd_bore_1_readen),
        .boreChildrenBd_bore_1_addr_rd(boreChildrenBd_bore_1_addr_rd),
        .boreChildrenBd_bore_1_outdata(boreChildrenBd_bore_1_outdata),
        .boreChildrenBd_bore_2_array(boreChildrenBd_bore_2_array),
        .boreChildrenBd_bore_2_all(boreChildrenBd_bore_2_all),
        .boreChildrenBd_bore_2_req(boreChildrenBd_bore_2_req),
        .boreChildrenBd_bore_2_ack(boreChildrenBd_bore_2_ack),
        .boreChildrenBd_bore_2_writeen(boreChildrenBd_bore_2_writeen),
        .boreChildrenBd_bore_2_be(boreChildrenBd_bore_2_be),
        .boreChildrenBd_bore_2_addr(boreChildrenBd_bore_2_addr),
        .boreChildrenBd_bore_2_indata(boreChildrenBd_bore_2_indata),
        .boreChildrenBd_bore_2_readen(boreChildrenBd_bore_2_readen),
        .boreChildrenBd_bore_2_addr_rd(boreChildrenBd_bore_2_addr_rd),
        .boreChildrenBd_bore_2_outdata(boreChildrenBd_bore_2_outdata),
        .boreChildrenBd_bore_3_array(boreChildrenBd_bore_3_array),
        .boreChildrenBd_bore_3_all(boreChildrenBd_bore_3_all),
        .boreChildrenBd_bore_3_req(boreChildrenBd_bore_3_req),
        .boreChildrenBd_bore_3_ack(boreChildrenBd_bore_3_ack),
        .boreChildrenBd_bore_3_writeen(boreChildrenBd_bore_3_writeen),
        .boreChildrenBd_bore_3_be(boreChildrenBd_bore_3_be),
        .boreChildrenBd_bore_3_addr(boreChildrenBd_bore_3_addr),
        .boreChildrenBd_bore_3_indata(boreChildrenBd_bore_3_indata),
        .boreChildrenBd_bore_3_readen(boreChildrenBd_bore_3_readen),
        .boreChildrenBd_bore_3_addr_rd(boreChildrenBd_bore_3_addr_rd),
        .boreChildrenBd_bore_3_outdata(boreChildrenBd_bore_3_outdata),
        .boreChildrenBd_bore_4_array(boreChildrenBd_bore_4_array),
        .boreChildrenBd_bore_4_all(boreChildrenBd_bore_4_all),
        .boreChildrenBd_bore_4_req(boreChildrenBd_bore_4_req),
        .boreChildrenBd_bore_4_ack(boreChildrenBd_bore_4_ack),
        .boreChildrenBd_bore_4_writeen(boreChildrenBd_bore_4_writeen),
        .boreChildrenBd_bore_4_be(boreChildrenBd_bore_4_be),
        .boreChildrenBd_bore_4_addr(boreChildrenBd_bore_4_addr),
        .boreChildrenBd_bore_4_indata(boreChildrenBd_bore_4_indata),
        .boreChildrenBd_bore_4_readen(boreChildrenBd_bore_4_readen),
        .boreChildrenBd_bore_4_addr_rd(boreChildrenBd_bore_4_addr_rd),
        .boreChildrenBd_bore_4_outdata(boreChildrenBd_bore_4_outdata),
        .boreChildrenBd_bore_5_addr(boreChildrenBd_bore_5_addr),
        .boreChildrenBd_bore_5_addr_rd(boreChildrenBd_bore_5_addr_rd),
        .boreChildrenBd_bore_5_wdata(boreChildrenBd_bore_5_wdata),
        .boreChildrenBd_bore_5_wmask(boreChildrenBd_bore_5_wmask),
        .boreChildrenBd_bore_5_re(boreChildrenBd_bore_5_re),
        .boreChildrenBd_bore_5_we(boreChildrenBd_bore_5_we),
        .boreChildrenBd_bore_5_rdata(boreChildrenBd_bore_5_rdata),
        .boreChildrenBd_bore_5_ack(boreChildrenBd_bore_5_ack),
        .boreChildrenBd_bore_5_selectedOH(boreChildrenBd_bore_5_selectedOH),
        .boreChildrenBd_bore_5_array(boreChildrenBd_bore_5_array),
        .boreChildrenBd_bore_6_addr(boreChildrenBd_bore_6_addr),
        .boreChildrenBd_bore_6_addr_rd(boreChildrenBd_bore_6_addr_rd),
        .boreChildrenBd_bore_6_wdata(boreChildrenBd_bore_6_wdata),
        .boreChildrenBd_bore_6_wmask(boreChildrenBd_bore_6_wmask),
        .boreChildrenBd_bore_6_re(boreChildrenBd_bore_6_re),
        .boreChildrenBd_bore_6_we(boreChildrenBd_bore_6_we),
        .boreChildrenBd_bore_6_rdata(boreChildrenBd_bore_6_rdata),
        .boreChildrenBd_bore_6_ack(boreChildrenBd_bore_6_ack),
        .boreChildrenBd_bore_6_selectedOH(boreChildrenBd_bore_6_selectedOH),
        .boreChildrenBd_bore_6_array(boreChildrenBd_bore_6_array),
        .boreChildrenBd_bore_7_addr(boreChildrenBd_bore_7_addr),
        .boreChildrenBd_bore_7_addr_rd(boreChildrenBd_bore_7_addr_rd),
        .boreChildrenBd_bore_7_wdata(boreChildrenBd_bore_7_wdata),
        .boreChildrenBd_bore_7_wmask(boreChildrenBd_bore_7_wmask),
        .boreChildrenBd_bore_7_re(boreChildrenBd_bore_7_re),
        .boreChildrenBd_bore_7_we(boreChildrenBd_bore_7_we),
        .boreChildrenBd_bore_7_rdata(boreChildrenBd_bore_7_rdata),
        .boreChildrenBd_bore_7_ack(boreChildrenBd_bore_7_ack),
        .boreChildrenBd_bore_7_selectedOH(boreChildrenBd_bore_7_selectedOH),
        .boreChildrenBd_bore_7_array(boreChildrenBd_bore_7_array),
        .boreChildrenBd_bore_8_addr(boreChildrenBd_bore_8_addr),
        .boreChildrenBd_bore_8_addr_rd(boreChildrenBd_bore_8_addr_rd),
        .boreChildrenBd_bore_8_wdata(boreChildrenBd_bore_8_wdata),
        .boreChildrenBd_bore_8_wmask(boreChildrenBd_bore_8_wmask),
        .boreChildrenBd_bore_8_re(boreChildrenBd_bore_8_re),
        .boreChildrenBd_bore_8_we(boreChildrenBd_bore_8_we),
        .boreChildrenBd_bore_8_rdata(boreChildrenBd_bore_8_rdata),
        .boreChildrenBd_bore_8_ack(boreChildrenBd_bore_8_ack),
        .boreChildrenBd_bore_8_selectedOH(boreChildrenBd_bore_8_selectedOH),
        .boreChildrenBd_bore_8_array(boreChildrenBd_bore_8_array),
        .boreChildrenBd_bore_9_addr(boreChildrenBd_bore_9_addr),
        .boreChildrenBd_bore_9_addr_rd(boreChildrenBd_bore_9_addr_rd),
        .boreChildrenBd_bore_9_wdata(boreChildrenBd_bore_9_wdata),
        .boreChildrenBd_bore_9_wmask(boreChildrenBd_bore_9_wmask),
        .boreChildrenBd_bore_9_re(boreChildrenBd_bore_9_re),
        .boreChildrenBd_bore_9_we(boreChildrenBd_bore_9_we),
        .boreChildrenBd_bore_9_rdata(boreChildrenBd_bore_9_rdata),
        .boreChildrenBd_bore_9_ack(boreChildrenBd_bore_9_ack),
        .boreChildrenBd_bore_9_selectedOH(boreChildrenBd_bore_9_selectedOH),
        .boreChildrenBd_bore_9_array(boreChildrenBd_bore_9_array),
        .boreChildrenBd_bore_10_addr(boreChildrenBd_bore_10_addr),
        .boreChildrenBd_bore_10_addr_rd(boreChildrenBd_bore_10_addr_rd),
        .boreChildrenBd_bore_10_wdata(boreChildrenBd_bore_10_wdata),
        .boreChildrenBd_bore_10_wmask(boreChildrenBd_bore_10_wmask),
        .boreChildrenBd_bore_10_re(boreChildrenBd_bore_10_re),
        .boreChildrenBd_bore_10_we(boreChildrenBd_bore_10_we),
        .boreChildrenBd_bore_10_rdata(boreChildrenBd_bore_10_rdata),
        .boreChildrenBd_bore_10_ack(boreChildrenBd_bore_10_ack),
        .boreChildrenBd_bore_10_selectedOH(boreChildrenBd_bore_10_selectedOH),
        .boreChildrenBd_bore_10_array(boreChildrenBd_bore_10_array),
        .boreChildrenBd_bore_11_addr(boreChildrenBd_bore_11_addr),
        .boreChildrenBd_bore_11_addr_rd(boreChildrenBd_bore_11_addr_rd),
        .boreChildrenBd_bore_11_wdata(boreChildrenBd_bore_11_wdata),
        .boreChildrenBd_bore_11_wmask(boreChildrenBd_bore_11_wmask),
        .boreChildrenBd_bore_11_re(boreChildrenBd_bore_11_re),
        .boreChildrenBd_bore_11_we(boreChildrenBd_bore_11_we),
        .boreChildrenBd_bore_11_rdata(boreChildrenBd_bore_11_rdata),
        .boreChildrenBd_bore_11_ack(boreChildrenBd_bore_11_ack),
        .boreChildrenBd_bore_11_selectedOH(boreChildrenBd_bore_11_selectedOH),
        .boreChildrenBd_bore_11_array(boreChildrenBd_bore_11_array),
        .boreChildrenBd_bore_12_addr(boreChildrenBd_bore_12_addr),
        .boreChildrenBd_bore_12_addr_rd(boreChildrenBd_bore_12_addr_rd),
        .boreChildrenBd_bore_12_wdata(boreChildrenBd_bore_12_wdata),
        .boreChildrenBd_bore_12_wmask(boreChildrenBd_bore_12_wmask),
        .boreChildrenBd_bore_12_re(boreChildrenBd_bore_12_re),
        .boreChildrenBd_bore_12_we(boreChildrenBd_bore_12_we),
        .boreChildrenBd_bore_12_rdata(boreChildrenBd_bore_12_rdata),
        .boreChildrenBd_bore_12_ack(boreChildrenBd_bore_12_ack),
        .boreChildrenBd_bore_12_selectedOH(boreChildrenBd_bore_12_selectedOH),
        .boreChildrenBd_bore_12_array(boreChildrenBd_bore_12_array),
        .boreChildrenBd_bore_13_addr(boreChildrenBd_bore_13_addr),
        .boreChildrenBd_bore_13_addr_rd(boreChildrenBd_bore_13_addr_rd),
        .boreChildrenBd_bore_13_wdata(boreChildrenBd_bore_13_wdata),
        .boreChildrenBd_bore_13_wmask(boreChildrenBd_bore_13_wmask),
        .boreChildrenBd_bore_13_re(boreChildrenBd_bore_13_re),
        .boreChildrenBd_bore_13_we(boreChildrenBd_bore_13_we),
        .boreChildrenBd_bore_13_rdata(boreChildrenBd_bore_13_rdata),
        .boreChildrenBd_bore_13_ack(boreChildrenBd_bore_13_ack),
        .boreChildrenBd_bore_13_selectedOH(boreChildrenBd_bore_13_selectedOH),
        .boreChildrenBd_bore_13_array(boreChildrenBd_bore_13_array),
        .boreChildrenBd_bore_14_addr(boreChildrenBd_bore_14_addr),
        .boreChildrenBd_bore_14_addr_rd(boreChildrenBd_bore_14_addr_rd),
        .boreChildrenBd_bore_14_wdata(boreChildrenBd_bore_14_wdata),
        .boreChildrenBd_bore_14_wmask(boreChildrenBd_bore_14_wmask),
        .boreChildrenBd_bore_14_re(boreChildrenBd_bore_14_re),
        .boreChildrenBd_bore_14_we(boreChildrenBd_bore_14_we),
        .boreChildrenBd_bore_14_rdata(boreChildrenBd_bore_14_rdata),
        .boreChildrenBd_bore_14_ack(boreChildrenBd_bore_14_ack),
        .boreChildrenBd_bore_14_selectedOH(boreChildrenBd_bore_14_selectedOH),
        .boreChildrenBd_bore_14_array(boreChildrenBd_bore_14_array),
        .boreChildrenBd_bore_15_addr(boreChildrenBd_bore_15_addr),
        .boreChildrenBd_bore_15_addr_rd(boreChildrenBd_bore_15_addr_rd),
        .boreChildrenBd_bore_15_wdata(boreChildrenBd_bore_15_wdata),
        .boreChildrenBd_bore_15_wmask(boreChildrenBd_bore_15_wmask),
        .boreChildrenBd_bore_15_re(boreChildrenBd_bore_15_re),
        .boreChildrenBd_bore_15_we(boreChildrenBd_bore_15_we),
        .boreChildrenBd_bore_15_rdata(boreChildrenBd_bore_15_rdata),
        .boreChildrenBd_bore_15_ack(boreChildrenBd_bore_15_ack),
        .boreChildrenBd_bore_15_selectedOH(boreChildrenBd_bore_15_selectedOH),
        .boreChildrenBd_bore_15_array(boreChildrenBd_bore_15_array),
        .boreChildrenBd_bore_16_addr(boreChildrenBd_bore_16_addr),
        .boreChildrenBd_bore_16_addr_rd(boreChildrenBd_bore_16_addr_rd),
        .boreChildrenBd_bore_16_wdata(boreChildrenBd_bore_16_wdata),
        .boreChildrenBd_bore_16_wmask(boreChildrenBd_bore_16_wmask),
        .boreChildrenBd_bore_16_re(boreChildrenBd_bore_16_re),
        .boreChildrenBd_bore_16_we(boreChildrenBd_bore_16_we),
        .boreChildrenBd_bore_16_rdata(boreChildrenBd_bore_16_rdata),
        .boreChildrenBd_bore_16_ack(boreChildrenBd_bore_16_ack),
        .boreChildrenBd_bore_16_selectedOH(boreChildrenBd_bore_16_selectedOH),
        .boreChildrenBd_bore_16_array(boreChildrenBd_bore_16_array),
        .boreChildrenBd_bore_17_addr(boreChildrenBd_bore_17_addr),
        .boreChildrenBd_bore_17_addr_rd(boreChildrenBd_bore_17_addr_rd),
        .boreChildrenBd_bore_17_wdata(boreChildrenBd_bore_17_wdata),
        .boreChildrenBd_bore_17_wmask(boreChildrenBd_bore_17_wmask),
        .boreChildrenBd_bore_17_re(boreChildrenBd_bore_17_re),
        .boreChildrenBd_bore_17_we(boreChildrenBd_bore_17_we),
        .boreChildrenBd_bore_17_rdata(boreChildrenBd_bore_17_rdata),
        .boreChildrenBd_bore_17_ack(boreChildrenBd_bore_17_ack),
        .boreChildrenBd_bore_17_selectedOH(boreChildrenBd_bore_17_selectedOH),
        .boreChildrenBd_bore_17_array(boreChildrenBd_bore_17_array),
        .boreChildrenBd_bore_18_addr(boreChildrenBd_bore_18_addr),
        .boreChildrenBd_bore_18_addr_rd(boreChildrenBd_bore_18_addr_rd),
        .boreChildrenBd_bore_18_wdata(boreChildrenBd_bore_18_wdata),
        .boreChildrenBd_bore_18_wmask(boreChildrenBd_bore_18_wmask),
        .boreChildrenBd_bore_18_re(boreChildrenBd_bore_18_re),
        .boreChildrenBd_bore_18_we(boreChildrenBd_bore_18_we),
        .boreChildrenBd_bore_18_rdata(boreChildrenBd_bore_18_rdata),
        .boreChildrenBd_bore_18_ack(boreChildrenBd_bore_18_ack),
        .boreChildrenBd_bore_18_selectedOH(boreChildrenBd_bore_18_selectedOH),
        .boreChildrenBd_bore_18_array(boreChildrenBd_bore_18_array),
        .sigFromSrams_bore_ram_hold(sigFromSrams_bore_ram_hold),
        .sigFromSrams_bore_ram_bypass(sigFromSrams_bore_ram_bypass),
        .sigFromSrams_bore_ram_bp_clken(sigFromSrams_bore_ram_bp_clken),
        .sigFromSrams_bore_ram_aux_clk(sigFromSrams_bore_ram_aux_clk),
        .sigFromSrams_bore_ram_aux_ckbp(sigFromSrams_bore_ram_aux_ckbp),
        .sigFromSrams_bore_ram_mcp_hold(sigFromSrams_bore_ram_mcp_hold),
        .sigFromSrams_bore_cgen(sigFromSrams_bore_cgen),
        .sigFromSrams_bore_1_ram_hold(sigFromSrams_bore_1_ram_hold),
        .sigFromSrams_bore_1_ram_bypass(sigFromSrams_bore_1_ram_bypass),
        .sigFromSrams_bore_1_ram_bp_clken(sigFromSrams_bore_1_ram_bp_clken),
        .sigFromSrams_bore_1_ram_aux_clk(sigFromSrams_bore_1_ram_aux_clk),
        .sigFromSrams_bore_1_ram_aux_ckbp(sigFromSrams_bore_1_ram_aux_ckbp),
        .sigFromSrams_bore_1_ram_mcp_hold(sigFromSrams_bore_1_ram_mcp_hold),
        .sigFromSrams_bore_1_cgen(sigFromSrams_bore_1_cgen),
        .sigFromSrams_bore_2_ram_hold(sigFromSrams_bore_2_ram_hold),
        .sigFromSrams_bore_2_ram_bypass(sigFromSrams_bore_2_ram_bypass),
        .sigFromSrams_bore_2_ram_bp_clken(sigFromSrams_bore_2_ram_bp_clken),
        .sigFromSrams_bore_2_ram_aux_clk(sigFromSrams_bore_2_ram_aux_clk),
        .sigFromSrams_bore_2_ram_aux_ckbp(sigFromSrams_bore_2_ram_aux_ckbp),
        .sigFromSrams_bore_2_ram_mcp_hold(sigFromSrams_bore_2_ram_mcp_hold),
        .sigFromSrams_bore_2_cgen(sigFromSrams_bore_2_cgen),
        .sigFromSrams_bore_3_ram_hold(sigFromSrams_bore_3_ram_hold),
        .sigFromSrams_bore_3_ram_bypass(sigFromSrams_bore_3_ram_bypass),
        .sigFromSrams_bore_3_ram_bp_clken(sigFromSrams_bore_3_ram_bp_clken),
        .sigFromSrams_bore_3_ram_aux_clk(sigFromSrams_bore_3_ram_aux_clk),
        .sigFromSrams_bore_3_ram_aux_ckbp(sigFromSrams_bore_3_ram_aux_ckbp),
        .sigFromSrams_bore_3_ram_mcp_hold(sigFromSrams_bore_3_ram_mcp_hold),
        .sigFromSrams_bore_3_cgen(sigFromSrams_bore_3_cgen),
        .sigFromSrams_bore_4_ram_hold(sigFromSrams_bore_4_ram_hold),
        .sigFromSrams_bore_4_ram_bypass(sigFromSrams_bore_4_ram_bypass),
        .sigFromSrams_bore_4_ram_bp_clken(sigFromSrams_bore_4_ram_bp_clken),
        .sigFromSrams_bore_4_ram_aux_clk(sigFromSrams_bore_4_ram_aux_clk),
        .sigFromSrams_bore_4_ram_aux_ckbp(sigFromSrams_bore_4_ram_aux_ckbp),
        .sigFromSrams_bore_4_ram_mcp_hold(sigFromSrams_bore_4_ram_mcp_hold),
        .sigFromSrams_bore_4_cgen(sigFromSrams_bore_4_cgen),
        .sigFromSrams_bore_5_ram_hold(sigFromSrams_bore_5_ram_hold),
        .sigFromSrams_bore_5_ram_bypass(sigFromSrams_bore_5_ram_bypass),
        .sigFromSrams_bore_5_ram_bp_clken(sigFromSrams_bore_5_ram_bp_clken),
        .sigFromSrams_bore_5_ram_aux_clk(sigFromSrams_bore_5_ram_aux_clk),
        .sigFromSrams_bore_5_ram_aux_ckbp(sigFromSrams_bore_5_ram_aux_ckbp),
        .sigFromSrams_bore_5_ram_mcp_hold(sigFromSrams_bore_5_ram_mcp_hold),
        .sigFromSrams_bore_5_cgen(sigFromSrams_bore_5_cgen),
        .sigFromSrams_bore_6_ram_hold(sigFromSrams_bore_6_ram_hold),
        .sigFromSrams_bore_6_ram_bypass(sigFromSrams_bore_6_ram_bypass),
        .sigFromSrams_bore_6_ram_bp_clken(sigFromSrams_bore_6_ram_bp_clken),
        .sigFromSrams_bore_6_ram_aux_clk(sigFromSrams_bore_6_ram_aux_clk),
        .sigFromSrams_bore_6_ram_aux_ckbp(sigFromSrams_bore_6_ram_aux_ckbp),
        .sigFromSrams_bore_6_ram_mcp_hold(sigFromSrams_bore_6_ram_mcp_hold),
        .sigFromSrams_bore_6_cgen(sigFromSrams_bore_6_cgen),
        .sigFromSrams_bore_7_ram_hold(sigFromSrams_bore_7_ram_hold),
        .sigFromSrams_bore_7_ram_bypass(sigFromSrams_bore_7_ram_bypass),
        .sigFromSrams_bore_7_ram_bp_clken(sigFromSrams_bore_7_ram_bp_clken),
        .sigFromSrams_bore_7_ram_aux_clk(sigFromSrams_bore_7_ram_aux_clk),
        .sigFromSrams_bore_7_ram_aux_ckbp(sigFromSrams_bore_7_ram_aux_ckbp),
        .sigFromSrams_bore_7_ram_mcp_hold(sigFromSrams_bore_7_ram_mcp_hold),
        .sigFromSrams_bore_7_cgen(sigFromSrams_bore_7_cgen),
        .sigFromSrams_bore_8_ram_hold(sigFromSrams_bore_8_ram_hold),
        .sigFromSrams_bore_8_ram_bypass(sigFromSrams_bore_8_ram_bypass),
        .sigFromSrams_bore_8_ram_bp_clken(sigFromSrams_bore_8_ram_bp_clken),
        .sigFromSrams_bore_8_ram_aux_clk(sigFromSrams_bore_8_ram_aux_clk),
        .sigFromSrams_bore_8_ram_aux_ckbp(sigFromSrams_bore_8_ram_aux_ckbp),
        .sigFromSrams_bore_8_ram_mcp_hold(sigFromSrams_bore_8_ram_mcp_hold),
        .sigFromSrams_bore_8_cgen(sigFromSrams_bore_8_cgen),
        .sigFromSrams_bore_9_ram_hold(sigFromSrams_bore_9_ram_hold),
        .sigFromSrams_bore_9_ram_bypass(sigFromSrams_bore_9_ram_bypass),
        .sigFromSrams_bore_9_ram_bp_clken(sigFromSrams_bore_9_ram_bp_clken),
        .sigFromSrams_bore_9_ram_aux_clk(sigFromSrams_bore_9_ram_aux_clk),
        .sigFromSrams_bore_9_ram_aux_ckbp(sigFromSrams_bore_9_ram_aux_ckbp),
        .sigFromSrams_bore_9_ram_mcp_hold(sigFromSrams_bore_9_ram_mcp_hold),
        .sigFromSrams_bore_9_cgen(sigFromSrams_bore_9_cgen),
        .sigFromSrams_bore_10_ram_hold(sigFromSrams_bore_10_ram_hold),
        .sigFromSrams_bore_10_ram_bypass(sigFromSrams_bore_10_ram_bypass),
        .sigFromSrams_bore_10_ram_bp_clken(sigFromSrams_bore_10_ram_bp_clken),
        .sigFromSrams_bore_10_ram_aux_clk(sigFromSrams_bore_10_ram_aux_clk),
        .sigFromSrams_bore_10_ram_aux_ckbp(sigFromSrams_bore_10_ram_aux_ckbp),
        .sigFromSrams_bore_10_ram_mcp_hold(sigFromSrams_bore_10_ram_mcp_hold),
        .sigFromSrams_bore_10_cgen(sigFromSrams_bore_10_cgen),
        .sigFromSrams_bore_11_ram_hold(sigFromSrams_bore_11_ram_hold),
        .sigFromSrams_bore_11_ram_bypass(sigFromSrams_bore_11_ram_bypass),
        .sigFromSrams_bore_11_ram_bp_clken(sigFromSrams_bore_11_ram_bp_clken),
        .sigFromSrams_bore_11_ram_aux_clk(sigFromSrams_bore_11_ram_aux_clk),
        .sigFromSrams_bore_11_ram_aux_ckbp(sigFromSrams_bore_11_ram_aux_ckbp),
        .sigFromSrams_bore_11_ram_mcp_hold(sigFromSrams_bore_11_ram_mcp_hold),
        .sigFromSrams_bore_11_cgen(sigFromSrams_bore_11_cgen),
        .sigFromSrams_bore_12_ram_hold(sigFromSrams_bore_12_ram_hold),
        .sigFromSrams_bore_12_ram_bypass(sigFromSrams_bore_12_ram_bypass),
        .sigFromSrams_bore_12_ram_bp_clken(sigFromSrams_bore_12_ram_bp_clken),
        .sigFromSrams_bore_12_ram_aux_clk(sigFromSrams_bore_12_ram_aux_clk),
        .sigFromSrams_bore_12_ram_aux_ckbp(sigFromSrams_bore_12_ram_aux_ckbp),
        .sigFromSrams_bore_12_ram_mcp_hold(sigFromSrams_bore_12_ram_mcp_hold),
        .sigFromSrams_bore_12_cgen(sigFromSrams_bore_12_cgen),
        .sigFromSrams_bore_13_ram_hold(sigFromSrams_bore_13_ram_hold),
        .sigFromSrams_bore_13_ram_bypass(sigFromSrams_bore_13_ram_bypass),
        .sigFromSrams_bore_13_ram_bp_clken(sigFromSrams_bore_13_ram_bp_clken),
        .sigFromSrams_bore_13_ram_aux_clk(sigFromSrams_bore_13_ram_aux_clk),
        .sigFromSrams_bore_13_ram_aux_ckbp(sigFromSrams_bore_13_ram_aux_ckbp),
        .sigFromSrams_bore_13_ram_mcp_hold(sigFromSrams_bore_13_ram_mcp_hold),
        .sigFromSrams_bore_13_cgen(sigFromSrams_bore_13_cgen),
        .sigFromSrams_bore_14_ram_hold(sigFromSrams_bore_14_ram_hold),
        .sigFromSrams_bore_14_ram_bypass(sigFromSrams_bore_14_ram_bypass),
        .sigFromSrams_bore_14_ram_bp_clken(sigFromSrams_bore_14_ram_bp_clken),
        .sigFromSrams_bore_14_ram_aux_clk(sigFromSrams_bore_14_ram_aux_clk),
        .sigFromSrams_bore_14_ram_aux_ckbp(sigFromSrams_bore_14_ram_aux_ckbp),
        .sigFromSrams_bore_14_ram_mcp_hold(sigFromSrams_bore_14_ram_mcp_hold),
        .sigFromSrams_bore_14_cgen(sigFromSrams_bore_14_cgen),
        .sigFromSrams_bore_15_ram_hold(sigFromSrams_bore_15_ram_hold),
        .sigFromSrams_bore_15_ram_bypass(sigFromSrams_bore_15_ram_bypass),
        .sigFromSrams_bore_15_ram_bp_clken(sigFromSrams_bore_15_ram_bp_clken),
        .sigFromSrams_bore_15_ram_aux_clk(sigFromSrams_bore_15_ram_aux_clk),
        .sigFromSrams_bore_15_ram_aux_ckbp(sigFromSrams_bore_15_ram_aux_ckbp),
        .sigFromSrams_bore_15_ram_mcp_hold(sigFromSrams_bore_15_ram_mcp_hold),
        .sigFromSrams_bore_15_cgen(sigFromSrams_bore_15_cgen),
        .sigFromSrams_bore_16_ram_hold(sigFromSrams_bore_16_ram_hold),
        .sigFromSrams_bore_16_ram_bypass(sigFromSrams_bore_16_ram_bypass),
        .sigFromSrams_bore_16_ram_bp_clken(sigFromSrams_bore_16_ram_bp_clken),
        .sigFromSrams_bore_16_ram_aux_clk(sigFromSrams_bore_16_ram_aux_clk),
        .sigFromSrams_bore_16_ram_aux_ckbp(sigFromSrams_bore_16_ram_aux_ckbp),
        .sigFromSrams_bore_16_ram_mcp_hold(sigFromSrams_bore_16_ram_mcp_hold),
        .sigFromSrams_bore_16_cgen(sigFromSrams_bore_16_cgen),
        .sigFromSrams_bore_17_ram_hold(sigFromSrams_bore_17_ram_hold),
        .sigFromSrams_bore_17_ram_bypass(sigFromSrams_bore_17_ram_bypass),
        .sigFromSrams_bore_17_ram_bp_clken(sigFromSrams_bore_17_ram_bp_clken),
        .sigFromSrams_bore_17_ram_aux_clk(sigFromSrams_bore_17_ram_aux_clk),
        .sigFromSrams_bore_17_ram_aux_ckbp(sigFromSrams_bore_17_ram_aux_ckbp),
        .sigFromSrams_bore_17_ram_mcp_hold(sigFromSrams_bore_17_ram_mcp_hold),
        .sigFromSrams_bore_17_cgen(sigFromSrams_bore_17_cgen),
        .sigFromSrams_bore_18_ram_hold(sigFromSrams_bore_18_ram_hold),
        .sigFromSrams_bore_18_ram_bypass(sigFromSrams_bore_18_ram_bypass),
        .sigFromSrams_bore_18_ram_bp_clken(sigFromSrams_bore_18_ram_bp_clken),
        .sigFromSrams_bore_18_ram_aux_clk(sigFromSrams_bore_18_ram_aux_clk),
        .sigFromSrams_bore_18_ram_aux_ckbp(sigFromSrams_bore_18_ram_aux_ckbp),
        .sigFromSrams_bore_18_ram_mcp_hold(sigFromSrams_bore_18_ram_mcp_hold),
        .sigFromSrams_bore_18_cgen(sigFromSrams_bore_18_cgen),
        .sigFromSrams_bore_19_ram_hold(sigFromSrams_bore_19_ram_hold),
        .sigFromSrams_bore_19_ram_bypass(sigFromSrams_bore_19_ram_bypass),
        .sigFromSrams_bore_19_ram_bp_clken(sigFromSrams_bore_19_ram_bp_clken),
        .sigFromSrams_bore_19_ram_aux_clk(sigFromSrams_bore_19_ram_aux_clk),
        .sigFromSrams_bore_19_ram_aux_ckbp(sigFromSrams_bore_19_ram_aux_ckbp),
        .sigFromSrams_bore_19_ram_mcp_hold(sigFromSrams_bore_19_ram_mcp_hold),
        .sigFromSrams_bore_19_cgen(sigFromSrams_bore_19_cgen),
        .sigFromSrams_bore_20_ram_hold(sigFromSrams_bore_20_ram_hold),
        .sigFromSrams_bore_20_ram_bypass(sigFromSrams_bore_20_ram_bypass),
        .sigFromSrams_bore_20_ram_bp_clken(sigFromSrams_bore_20_ram_bp_clken),
        .sigFromSrams_bore_20_ram_aux_clk(sigFromSrams_bore_20_ram_aux_clk),
        .sigFromSrams_bore_20_ram_aux_ckbp(sigFromSrams_bore_20_ram_aux_ckbp),
        .sigFromSrams_bore_20_ram_mcp_hold(sigFromSrams_bore_20_ram_mcp_hold),
        .sigFromSrams_bore_20_cgen(sigFromSrams_bore_20_cgen),
        .sigFromSrams_bore_21_ram_hold(sigFromSrams_bore_21_ram_hold),
        .sigFromSrams_bore_21_ram_bypass(sigFromSrams_bore_21_ram_bypass),
        .sigFromSrams_bore_21_ram_bp_clken(sigFromSrams_bore_21_ram_bp_clken),
        .sigFromSrams_bore_21_ram_aux_clk(sigFromSrams_bore_21_ram_aux_clk),
        .sigFromSrams_bore_21_ram_aux_ckbp(sigFromSrams_bore_21_ram_aux_ckbp),
        .sigFromSrams_bore_21_ram_mcp_hold(sigFromSrams_bore_21_ram_mcp_hold),
        .sigFromSrams_bore_21_cgen(sigFromSrams_bore_21_cgen),
        .sigFromSrams_bore_22_ram_hold(sigFromSrams_bore_22_ram_hold),
        .sigFromSrams_bore_22_ram_bypass(sigFromSrams_bore_22_ram_bypass),
        .sigFromSrams_bore_22_ram_bp_clken(sigFromSrams_bore_22_ram_bp_clken),
        .sigFromSrams_bore_22_ram_aux_clk(sigFromSrams_bore_22_ram_aux_clk),
        .sigFromSrams_bore_22_ram_aux_ckbp(sigFromSrams_bore_22_ram_aux_ckbp),
        .sigFromSrams_bore_22_ram_mcp_hold(sigFromSrams_bore_22_ram_mcp_hold),
        .sigFromSrams_bore_22_cgen(sigFromSrams_bore_22_cgen),
        .sigFromSrams_bore_23_ram_hold(sigFromSrams_bore_23_ram_hold),
        .sigFromSrams_bore_23_ram_bypass(sigFromSrams_bore_23_ram_bypass),
        .sigFromSrams_bore_23_ram_bp_clken(sigFromSrams_bore_23_ram_bp_clken),
        .sigFromSrams_bore_23_ram_aux_clk(sigFromSrams_bore_23_ram_aux_clk),
        .sigFromSrams_bore_23_ram_aux_ckbp(sigFromSrams_bore_23_ram_aux_ckbp),
        .sigFromSrams_bore_23_ram_mcp_hold(sigFromSrams_bore_23_ram_mcp_hold),
        .sigFromSrams_bore_23_cgen(sigFromSrams_bore_23_cgen),
        .sigFromSrams_bore_24_ram_hold(sigFromSrams_bore_24_ram_hold),
        .sigFromSrams_bore_24_ram_bypass(sigFromSrams_bore_24_ram_bypass),
        .sigFromSrams_bore_24_ram_bp_clken(sigFromSrams_bore_24_ram_bp_clken),
        .sigFromSrams_bore_24_ram_aux_clk(sigFromSrams_bore_24_ram_aux_clk),
        .sigFromSrams_bore_24_ram_aux_ckbp(sigFromSrams_bore_24_ram_aux_ckbp),
        .sigFromSrams_bore_24_ram_mcp_hold(sigFromSrams_bore_24_ram_mcp_hold),
        .sigFromSrams_bore_24_cgen(sigFromSrams_bore_24_cgen),
        .sigFromSrams_bore_25_ram_hold(sigFromSrams_bore_25_ram_hold),
        .sigFromSrams_bore_25_ram_bypass(sigFromSrams_bore_25_ram_bypass),
        .sigFromSrams_bore_25_ram_bp_clken(sigFromSrams_bore_25_ram_bp_clken),
        .sigFromSrams_bore_25_ram_aux_clk(sigFromSrams_bore_25_ram_aux_clk),
        .sigFromSrams_bore_25_ram_aux_ckbp(sigFromSrams_bore_25_ram_aux_ckbp),
        .sigFromSrams_bore_25_ram_mcp_hold(sigFromSrams_bore_25_ram_mcp_hold),
        .sigFromSrams_bore_25_cgen(sigFromSrams_bore_25_cgen),
        .sigFromSrams_bore_26_ram_hold(sigFromSrams_bore_26_ram_hold),
        .sigFromSrams_bore_26_ram_bypass(sigFromSrams_bore_26_ram_bypass),
        .sigFromSrams_bore_26_ram_bp_clken(sigFromSrams_bore_26_ram_bp_clken),
        .sigFromSrams_bore_26_ram_aux_clk(sigFromSrams_bore_26_ram_aux_clk),
        .sigFromSrams_bore_26_ram_aux_ckbp(sigFromSrams_bore_26_ram_aux_ckbp),
        .sigFromSrams_bore_26_ram_mcp_hold(sigFromSrams_bore_26_ram_mcp_hold),
        .sigFromSrams_bore_26_cgen(sigFromSrams_bore_26_cgen),
        .sigFromSrams_bore_27_ram_hold(sigFromSrams_bore_27_ram_hold),
        .sigFromSrams_bore_27_ram_bypass(sigFromSrams_bore_27_ram_bypass),
        .sigFromSrams_bore_27_ram_bp_clken(sigFromSrams_bore_27_ram_bp_clken),
        .sigFromSrams_bore_27_ram_aux_clk(sigFromSrams_bore_27_ram_aux_clk),
        .sigFromSrams_bore_27_ram_aux_ckbp(sigFromSrams_bore_27_ram_aux_ckbp),
        .sigFromSrams_bore_27_ram_mcp_hold(sigFromSrams_bore_27_ram_mcp_hold),
        .sigFromSrams_bore_27_cgen(sigFromSrams_bore_27_cgen),
        .sigFromSrams_bore_28_ram_hold(sigFromSrams_bore_28_ram_hold),
        .sigFromSrams_bore_28_ram_bypass(sigFromSrams_bore_28_ram_bypass),
        .sigFromSrams_bore_28_ram_bp_clken(sigFromSrams_bore_28_ram_bp_clken),
        .sigFromSrams_bore_28_ram_aux_clk(sigFromSrams_bore_28_ram_aux_clk),
        .sigFromSrams_bore_28_ram_aux_ckbp(sigFromSrams_bore_28_ram_aux_ckbp),
        .sigFromSrams_bore_28_ram_mcp_hold(sigFromSrams_bore_28_ram_mcp_hold),
        .sigFromSrams_bore_28_cgen(sigFromSrams_bore_28_cgen),
        .sigFromSrams_bore_29_ram_hold(sigFromSrams_bore_29_ram_hold),
        .sigFromSrams_bore_29_ram_bypass(sigFromSrams_bore_29_ram_bypass),
        .sigFromSrams_bore_29_ram_bp_clken(sigFromSrams_bore_29_ram_bp_clken),
        .sigFromSrams_bore_29_ram_aux_clk(sigFromSrams_bore_29_ram_aux_clk),
        .sigFromSrams_bore_29_ram_aux_ckbp(sigFromSrams_bore_29_ram_aux_ckbp),
        .sigFromSrams_bore_29_ram_mcp_hold(sigFromSrams_bore_29_ram_mcp_hold),
        .sigFromSrams_bore_29_cgen(sigFromSrams_bore_29_cgen),
        .sigFromSrams_bore_30_ram_hold(sigFromSrams_bore_30_ram_hold),
        .sigFromSrams_bore_30_ram_bypass(sigFromSrams_bore_30_ram_bypass),
        .sigFromSrams_bore_30_ram_bp_clken(sigFromSrams_bore_30_ram_bp_clken),
        .sigFromSrams_bore_30_ram_aux_clk(sigFromSrams_bore_30_ram_aux_clk),
        .sigFromSrams_bore_30_ram_aux_ckbp(sigFromSrams_bore_30_ram_aux_ckbp),
        .sigFromSrams_bore_30_ram_mcp_hold(sigFromSrams_bore_30_ram_mcp_hold),
        .sigFromSrams_bore_30_cgen(sigFromSrams_bore_30_cgen),
        .sigFromSrams_bore_31_ram_hold(sigFromSrams_bore_31_ram_hold),
        .sigFromSrams_bore_31_ram_bypass(sigFromSrams_bore_31_ram_bypass),
        .sigFromSrams_bore_31_ram_bp_clken(sigFromSrams_bore_31_ram_bp_clken),
        .sigFromSrams_bore_31_ram_aux_clk(sigFromSrams_bore_31_ram_aux_clk),
        .sigFromSrams_bore_31_ram_aux_ckbp(sigFromSrams_bore_31_ram_aux_ckbp),
        .sigFromSrams_bore_31_ram_mcp_hold(sigFromSrams_bore_31_ram_mcp_hold),
        .sigFromSrams_bore_31_cgen(sigFromSrams_bore_31_cgen),
        .sigFromSrams_bore_32_ram_hold(sigFromSrams_bore_32_ram_hold),
        .sigFromSrams_bore_32_ram_bypass(sigFromSrams_bore_32_ram_bypass),
        .sigFromSrams_bore_32_ram_bp_clken(sigFromSrams_bore_32_ram_bp_clken),
        .sigFromSrams_bore_32_ram_aux_clk(sigFromSrams_bore_32_ram_aux_clk),
        .sigFromSrams_bore_32_ram_aux_ckbp(sigFromSrams_bore_32_ram_aux_ckbp),
        .sigFromSrams_bore_32_ram_mcp_hold(sigFromSrams_bore_32_ram_mcp_hold),
        .sigFromSrams_bore_32_cgen(sigFromSrams_bore_32_cgen),
        .sigFromSrams_bore_33_ram_hold(sigFromSrams_bore_33_ram_hold),
        .sigFromSrams_bore_33_ram_bypass(sigFromSrams_bore_33_ram_bypass),
        .sigFromSrams_bore_33_ram_bp_clken(sigFromSrams_bore_33_ram_bp_clken),
        .sigFromSrams_bore_33_ram_aux_clk(sigFromSrams_bore_33_ram_aux_clk),
        .sigFromSrams_bore_33_ram_aux_ckbp(sigFromSrams_bore_33_ram_aux_ckbp),
        .sigFromSrams_bore_33_ram_mcp_hold(sigFromSrams_bore_33_ram_mcp_hold),
        .sigFromSrams_bore_33_cgen(sigFromSrams_bore_33_cgen),
        .sigFromSrams_bore_34_ram_hold(sigFromSrams_bore_34_ram_hold),
        .sigFromSrams_bore_34_ram_bypass(sigFromSrams_bore_34_ram_bypass),
        .sigFromSrams_bore_34_ram_bp_clken(sigFromSrams_bore_34_ram_bp_clken),
        .sigFromSrams_bore_34_ram_aux_clk(sigFromSrams_bore_34_ram_aux_clk),
        .sigFromSrams_bore_34_ram_aux_ckbp(sigFromSrams_bore_34_ram_aux_ckbp),
        .sigFromSrams_bore_34_ram_mcp_hold(sigFromSrams_bore_34_ram_mcp_hold),
        .sigFromSrams_bore_34_cgen(sigFromSrams_bore_34_cgen),
        .sigFromSrams_bore_35_ram_hold(sigFromSrams_bore_35_ram_hold),
        .sigFromSrams_bore_35_ram_bypass(sigFromSrams_bore_35_ram_bypass),
        .sigFromSrams_bore_35_ram_bp_clken(sigFromSrams_bore_35_ram_bp_clken),
        .sigFromSrams_bore_35_ram_aux_clk(sigFromSrams_bore_35_ram_aux_clk),
        .sigFromSrams_bore_35_ram_aux_ckbp(sigFromSrams_bore_35_ram_aux_ckbp),
        .sigFromSrams_bore_35_ram_mcp_hold(sigFromSrams_bore_35_ram_mcp_hold),
        .sigFromSrams_bore_35_cgen(sigFromSrams_bore_35_cgen),
        .sigFromSrams_bore_36_ram_hold(sigFromSrams_bore_36_ram_hold),
        .sigFromSrams_bore_36_ram_bypass(sigFromSrams_bore_36_ram_bypass),
        .sigFromSrams_bore_36_ram_bp_clken(sigFromSrams_bore_36_ram_bp_clken),
        .sigFromSrams_bore_36_ram_aux_clk(sigFromSrams_bore_36_ram_aux_clk),
        .sigFromSrams_bore_36_ram_aux_ckbp(sigFromSrams_bore_36_ram_aux_ckbp),
        .sigFromSrams_bore_36_ram_mcp_hold(sigFromSrams_bore_36_ram_mcp_hold),
        .sigFromSrams_bore_36_cgen(sigFromSrams_bore_36_cgen),
        .sigFromSrams_bore_37_ram_hold(sigFromSrams_bore_37_ram_hold),
        .sigFromSrams_bore_37_ram_bypass(sigFromSrams_bore_37_ram_bypass),
        .sigFromSrams_bore_37_ram_bp_clken(sigFromSrams_bore_37_ram_bp_clken),
        .sigFromSrams_bore_37_ram_aux_clk(sigFromSrams_bore_37_ram_aux_clk),
        .sigFromSrams_bore_37_ram_aux_ckbp(sigFromSrams_bore_37_ram_aux_ckbp),
        .sigFromSrams_bore_37_ram_mcp_hold(sigFromSrams_bore_37_ram_mcp_hold),
        .sigFromSrams_bore_37_cgen(sigFromSrams_bore_37_cgen),
        .sigFromSrams_bore_38_ram_hold(sigFromSrams_bore_38_ram_hold),
        .sigFromSrams_bore_38_ram_bypass(sigFromSrams_bore_38_ram_bypass),
        .sigFromSrams_bore_38_ram_bp_clken(sigFromSrams_bore_38_ram_bp_clken),
        .sigFromSrams_bore_38_ram_aux_clk(sigFromSrams_bore_38_ram_aux_clk),
        .sigFromSrams_bore_38_ram_aux_ckbp(sigFromSrams_bore_38_ram_aux_ckbp),
        .sigFromSrams_bore_38_ram_mcp_hold(sigFromSrams_bore_38_ram_mcp_hold),
        .sigFromSrams_bore_38_cgen(sigFromSrams_bore_38_cgen),
        .sigFromSrams_bore_39_ram_hold(sigFromSrams_bore_39_ram_hold),
        .sigFromSrams_bore_39_ram_bypass(sigFromSrams_bore_39_ram_bypass),
        .sigFromSrams_bore_39_ram_bp_clken(sigFromSrams_bore_39_ram_bp_clken),
        .sigFromSrams_bore_39_ram_aux_clk(sigFromSrams_bore_39_ram_aux_clk),
        .sigFromSrams_bore_39_ram_aux_ckbp(sigFromSrams_bore_39_ram_aux_ckbp),
        .sigFromSrams_bore_39_ram_mcp_hold(sigFromSrams_bore_39_ram_mcp_hold),
        .sigFromSrams_bore_39_cgen(sigFromSrams_bore_39_cgen),
        .sigFromSrams_bore_40_ram_hold(sigFromSrams_bore_40_ram_hold),
        .sigFromSrams_bore_40_ram_bypass(sigFromSrams_bore_40_ram_bypass),
        .sigFromSrams_bore_40_ram_bp_clken(sigFromSrams_bore_40_ram_bp_clken),
        .sigFromSrams_bore_40_ram_aux_clk(sigFromSrams_bore_40_ram_aux_clk),
        .sigFromSrams_bore_40_ram_aux_ckbp(sigFromSrams_bore_40_ram_aux_ckbp),
        .sigFromSrams_bore_40_ram_mcp_hold(sigFromSrams_bore_40_ram_mcp_hold),
        .sigFromSrams_bore_40_cgen(sigFromSrams_bore_40_cgen),
        .sigFromSrams_bore_41_ram_hold(sigFromSrams_bore_41_ram_hold),
        .sigFromSrams_bore_41_ram_bypass(sigFromSrams_bore_41_ram_bypass),
        .sigFromSrams_bore_41_ram_bp_clken(sigFromSrams_bore_41_ram_bp_clken),
        .sigFromSrams_bore_41_ram_aux_clk(sigFromSrams_bore_41_ram_aux_clk),
        .sigFromSrams_bore_41_ram_aux_ckbp(sigFromSrams_bore_41_ram_aux_ckbp),
        .sigFromSrams_bore_41_ram_mcp_hold(sigFromSrams_bore_41_ram_mcp_hold),
        .sigFromSrams_bore_41_cgen(sigFromSrams_bore_41_cgen),
        .sigFromSrams_bore_42_ram_hold(sigFromSrams_bore_42_ram_hold),
        .sigFromSrams_bore_42_ram_bypass(sigFromSrams_bore_42_ram_bypass),
        .sigFromSrams_bore_42_ram_bp_clken(sigFromSrams_bore_42_ram_bp_clken),
        .sigFromSrams_bore_42_ram_aux_clk(sigFromSrams_bore_42_ram_aux_clk),
        .sigFromSrams_bore_42_ram_aux_ckbp(sigFromSrams_bore_42_ram_aux_ckbp),
        .sigFromSrams_bore_42_ram_mcp_hold(sigFromSrams_bore_42_ram_mcp_hold),
        .sigFromSrams_bore_42_cgen(sigFromSrams_bore_42_cgen),
        .sigFromSrams_bore_43_ram_hold(sigFromSrams_bore_43_ram_hold),
        .sigFromSrams_bore_43_ram_bypass(sigFromSrams_bore_43_ram_bypass),
        .sigFromSrams_bore_43_ram_bp_clken(sigFromSrams_bore_43_ram_bp_clken),
        .sigFromSrams_bore_43_ram_aux_clk(sigFromSrams_bore_43_ram_aux_clk),
        .sigFromSrams_bore_43_ram_aux_ckbp(sigFromSrams_bore_43_ram_aux_ckbp),
        .sigFromSrams_bore_43_ram_mcp_hold(sigFromSrams_bore_43_ram_mcp_hold),
        .sigFromSrams_bore_43_cgen(sigFromSrams_bore_43_cgen),
        .sigFromSrams_bore_44_ram_hold(sigFromSrams_bore_44_ram_hold),
        .sigFromSrams_bore_44_ram_bypass(sigFromSrams_bore_44_ram_bypass),
        .sigFromSrams_bore_44_ram_bp_clken(sigFromSrams_bore_44_ram_bp_clken),
        .sigFromSrams_bore_44_ram_aux_clk(sigFromSrams_bore_44_ram_aux_clk),
        .sigFromSrams_bore_44_ram_aux_ckbp(sigFromSrams_bore_44_ram_aux_ckbp),
        .sigFromSrams_bore_44_ram_mcp_hold(sigFromSrams_bore_44_ram_mcp_hold),
        .sigFromSrams_bore_44_cgen(sigFromSrams_bore_44_cgen),
        .sigFromSrams_bore_45_ram_hold(sigFromSrams_bore_45_ram_hold),
        .sigFromSrams_bore_45_ram_bypass(sigFromSrams_bore_45_ram_bypass),
        .sigFromSrams_bore_45_ram_bp_clken(sigFromSrams_bore_45_ram_bp_clken),
        .sigFromSrams_bore_45_ram_aux_clk(sigFromSrams_bore_45_ram_aux_clk),
        .sigFromSrams_bore_45_ram_aux_ckbp(sigFromSrams_bore_45_ram_aux_ckbp),
        .sigFromSrams_bore_45_ram_mcp_hold(sigFromSrams_bore_45_ram_mcp_hold),
        .sigFromSrams_bore_45_cgen(sigFromSrams_bore_45_cgen),
        .sigFromSrams_bore_46_ram_hold(sigFromSrams_bore_46_ram_hold),
        .sigFromSrams_bore_46_ram_bypass(sigFromSrams_bore_46_ram_bypass),
        .sigFromSrams_bore_46_ram_bp_clken(sigFromSrams_bore_46_ram_bp_clken),
        .sigFromSrams_bore_46_ram_aux_clk(sigFromSrams_bore_46_ram_aux_clk),
        .sigFromSrams_bore_46_ram_aux_ckbp(sigFromSrams_bore_46_ram_aux_ckbp),
        .sigFromSrams_bore_46_ram_mcp_hold(sigFromSrams_bore_46_ram_mcp_hold),
        .sigFromSrams_bore_46_cgen(sigFromSrams_bore_46_cgen),
        .sigFromSrams_bore_47_ram_hold(sigFromSrams_bore_47_ram_hold),
        .sigFromSrams_bore_47_ram_bypass(sigFromSrams_bore_47_ram_bypass),
        .sigFromSrams_bore_47_ram_bp_clken(sigFromSrams_bore_47_ram_bp_clken),
        .sigFromSrams_bore_47_ram_aux_clk(sigFromSrams_bore_47_ram_aux_clk),
        .sigFromSrams_bore_47_ram_aux_ckbp(sigFromSrams_bore_47_ram_aux_ckbp),
        .sigFromSrams_bore_47_ram_mcp_hold(sigFromSrams_bore_47_ram_mcp_hold),
        .sigFromSrams_bore_47_cgen(sigFromSrams_bore_47_cgen),
        .sigFromSrams_bore_48_ram_hold(sigFromSrams_bore_48_ram_hold),
        .sigFromSrams_bore_48_ram_bypass(sigFromSrams_bore_48_ram_bypass),
        .sigFromSrams_bore_48_ram_bp_clken(sigFromSrams_bore_48_ram_bp_clken),
        .sigFromSrams_bore_48_ram_aux_clk(sigFromSrams_bore_48_ram_aux_clk),
        .sigFromSrams_bore_48_ram_aux_ckbp(sigFromSrams_bore_48_ram_aux_ckbp),
        .sigFromSrams_bore_48_ram_mcp_hold(sigFromSrams_bore_48_ram_mcp_hold),
        .sigFromSrams_bore_48_cgen(sigFromSrams_bore_48_cgen),
        .sigFromSrams_bore_49_ram_hold(sigFromSrams_bore_49_ram_hold),
        .sigFromSrams_bore_49_ram_bypass(sigFromSrams_bore_49_ram_bypass),
        .sigFromSrams_bore_49_ram_bp_clken(sigFromSrams_bore_49_ram_bp_clken),
        .sigFromSrams_bore_49_ram_aux_clk(sigFromSrams_bore_49_ram_aux_clk),
        .sigFromSrams_bore_49_ram_aux_ckbp(sigFromSrams_bore_49_ram_aux_ckbp),
        .sigFromSrams_bore_49_ram_mcp_hold(sigFromSrams_bore_49_ram_mcp_hold),
        .sigFromSrams_bore_49_cgen(sigFromSrams_bore_49_cgen),
        .sigFromSrams_bore_50_ram_hold(sigFromSrams_bore_50_ram_hold),
        .sigFromSrams_bore_50_ram_bypass(sigFromSrams_bore_50_ram_bypass),
        .sigFromSrams_bore_50_ram_bp_clken(sigFromSrams_bore_50_ram_bp_clken),
        .sigFromSrams_bore_50_ram_aux_clk(sigFromSrams_bore_50_ram_aux_clk),
        .sigFromSrams_bore_50_ram_aux_ckbp(sigFromSrams_bore_50_ram_aux_ckbp),
        .sigFromSrams_bore_50_ram_mcp_hold(sigFromSrams_bore_50_ram_mcp_hold),
        .sigFromSrams_bore_50_cgen(sigFromSrams_bore_50_cgen),
        .sigFromSrams_bore_51_ram_hold(sigFromSrams_bore_51_ram_hold),
        .sigFromSrams_bore_51_ram_bypass(sigFromSrams_bore_51_ram_bypass),
        .sigFromSrams_bore_51_ram_bp_clken(sigFromSrams_bore_51_ram_bp_clken),
        .sigFromSrams_bore_51_ram_aux_clk(sigFromSrams_bore_51_ram_aux_clk),
        .sigFromSrams_bore_51_ram_aux_ckbp(sigFromSrams_bore_51_ram_aux_ckbp),
        .sigFromSrams_bore_51_ram_mcp_hold(sigFromSrams_bore_51_ram_mcp_hold),
        .sigFromSrams_bore_51_cgen(sigFromSrams_bore_51_cgen),
        .sigFromSrams_bore_52_ram_hold(sigFromSrams_bore_52_ram_hold),
        .sigFromSrams_bore_52_ram_bypass(sigFromSrams_bore_52_ram_bypass),
        .sigFromSrams_bore_52_ram_bp_clken(sigFromSrams_bore_52_ram_bp_clken),
        .sigFromSrams_bore_52_ram_aux_clk(sigFromSrams_bore_52_ram_aux_clk),
        .sigFromSrams_bore_52_ram_aux_ckbp(sigFromSrams_bore_52_ram_aux_ckbp),
        .sigFromSrams_bore_52_ram_mcp_hold(sigFromSrams_bore_52_ram_mcp_hold),
        .sigFromSrams_bore_52_cgen(sigFromSrams_bore_52_cgen),
        .sigFromSrams_bore_53_ram_hold(sigFromSrams_bore_53_ram_hold),
        .sigFromSrams_bore_53_ram_bypass(sigFromSrams_bore_53_ram_bypass),
        .sigFromSrams_bore_53_ram_bp_clken(sigFromSrams_bore_53_ram_bp_clken),
        .sigFromSrams_bore_53_ram_aux_clk(sigFromSrams_bore_53_ram_aux_clk),
        .sigFromSrams_bore_53_ram_aux_ckbp(sigFromSrams_bore_53_ram_aux_ckbp),
        .sigFromSrams_bore_53_ram_mcp_hold(sigFromSrams_bore_53_ram_mcp_hold),
        .sigFromSrams_bore_53_cgen(sigFromSrams_bore_53_cgen),
        .sigFromSrams_bore_54_ram_hold(sigFromSrams_bore_54_ram_hold),
        .sigFromSrams_bore_54_ram_bypass(sigFromSrams_bore_54_ram_bypass),
        .sigFromSrams_bore_54_ram_bp_clken(sigFromSrams_bore_54_ram_bp_clken),
        .sigFromSrams_bore_54_ram_aux_clk(sigFromSrams_bore_54_ram_aux_clk),
        .sigFromSrams_bore_54_ram_aux_ckbp(sigFromSrams_bore_54_ram_aux_ckbp),
        .sigFromSrams_bore_54_ram_mcp_hold(sigFromSrams_bore_54_ram_mcp_hold),
        .sigFromSrams_bore_54_cgen(sigFromSrams_bore_54_cgen),
        .sigFromSrams_bore_55_ram_hold(sigFromSrams_bore_55_ram_hold),
        .sigFromSrams_bore_55_ram_bypass(sigFromSrams_bore_55_ram_bypass),
        .sigFromSrams_bore_55_ram_bp_clken(sigFromSrams_bore_55_ram_bp_clken),
        .sigFromSrams_bore_55_ram_aux_clk(sigFromSrams_bore_55_ram_aux_clk),
        .sigFromSrams_bore_55_ram_aux_ckbp(sigFromSrams_bore_55_ram_aux_ckbp),
        .sigFromSrams_bore_55_ram_mcp_hold(sigFromSrams_bore_55_ram_mcp_hold),
        .sigFromSrams_bore_55_cgen(sigFromSrams_bore_55_cgen),
        .sigFromSrams_bore_56_ram_hold(sigFromSrams_bore_56_ram_hold),
        .sigFromSrams_bore_56_ram_bypass(sigFromSrams_bore_56_ram_bypass),
        .sigFromSrams_bore_56_ram_bp_clken(sigFromSrams_bore_56_ram_bp_clken),
        .sigFromSrams_bore_56_ram_aux_clk(sigFromSrams_bore_56_ram_aux_clk),
        .sigFromSrams_bore_56_ram_aux_ckbp(sigFromSrams_bore_56_ram_aux_ckbp),
        .sigFromSrams_bore_56_ram_mcp_hold(sigFromSrams_bore_56_ram_mcp_hold),
        .sigFromSrams_bore_56_cgen(sigFromSrams_bore_56_cgen),
        .sigFromSrams_bore_57_ram_hold(sigFromSrams_bore_57_ram_hold),
        .sigFromSrams_bore_57_ram_bypass(sigFromSrams_bore_57_ram_bypass),
        .sigFromSrams_bore_57_ram_bp_clken(sigFromSrams_bore_57_ram_bp_clken),
        .sigFromSrams_bore_57_ram_aux_clk(sigFromSrams_bore_57_ram_aux_clk),
        .sigFromSrams_bore_57_ram_aux_ckbp(sigFromSrams_bore_57_ram_aux_ckbp),
        .sigFromSrams_bore_57_ram_mcp_hold(sigFromSrams_bore_57_ram_mcp_hold),
        .sigFromSrams_bore_57_cgen(sigFromSrams_bore_57_cgen),
        .sigFromSrams_bore_58_ram_hold(sigFromSrams_bore_58_ram_hold),
        .sigFromSrams_bore_58_ram_bypass(sigFromSrams_bore_58_ram_bypass),
        .sigFromSrams_bore_58_ram_bp_clken(sigFromSrams_bore_58_ram_bp_clken),
        .sigFromSrams_bore_58_ram_aux_clk(sigFromSrams_bore_58_ram_aux_clk),
        .sigFromSrams_bore_58_ram_aux_ckbp(sigFromSrams_bore_58_ram_aux_ckbp),
        .sigFromSrams_bore_58_ram_mcp_hold(sigFromSrams_bore_58_ram_mcp_hold),
        .sigFromSrams_bore_58_cgen(sigFromSrams_bore_58_cgen),
        .sigFromSrams_bore_59_ram_hold(sigFromSrams_bore_59_ram_hold),
        .sigFromSrams_bore_59_ram_bypass(sigFromSrams_bore_59_ram_bypass),
        .sigFromSrams_bore_59_ram_bp_clken(sigFromSrams_bore_59_ram_bp_clken),
        .sigFromSrams_bore_59_ram_aux_clk(sigFromSrams_bore_59_ram_aux_clk),
        .sigFromSrams_bore_59_ram_aux_ckbp(sigFromSrams_bore_59_ram_aux_ckbp),
        .sigFromSrams_bore_59_ram_mcp_hold(sigFromSrams_bore_59_ram_mcp_hold),
        .sigFromSrams_bore_59_cgen(sigFromSrams_bore_59_cgen),
        .sigFromSrams_bore_60_ram_hold(sigFromSrams_bore_60_ram_hold),
        .sigFromSrams_bore_60_ram_bypass(sigFromSrams_bore_60_ram_bypass),
        .sigFromSrams_bore_60_ram_bp_clken(sigFromSrams_bore_60_ram_bp_clken),
        .sigFromSrams_bore_60_ram_aux_clk(sigFromSrams_bore_60_ram_aux_clk),
        .sigFromSrams_bore_60_ram_aux_ckbp(sigFromSrams_bore_60_ram_aux_ckbp),
        .sigFromSrams_bore_60_ram_mcp_hold(sigFromSrams_bore_60_ram_mcp_hold),
        .sigFromSrams_bore_60_cgen(sigFromSrams_bore_60_cgen),
        .sigFromSrams_bore_61_ram_hold(sigFromSrams_bore_61_ram_hold),
        .sigFromSrams_bore_61_ram_bypass(sigFromSrams_bore_61_ram_bypass),
        .sigFromSrams_bore_61_ram_bp_clken(sigFromSrams_bore_61_ram_bp_clken),
        .sigFromSrams_bore_61_ram_aux_clk(sigFromSrams_bore_61_ram_aux_clk),
        .sigFromSrams_bore_61_ram_aux_ckbp(sigFromSrams_bore_61_ram_aux_ckbp),
        .sigFromSrams_bore_61_ram_mcp_hold(sigFromSrams_bore_61_ram_mcp_hold),
        .sigFromSrams_bore_61_cgen(sigFromSrams_bore_61_cgen),
        .sigFromSrams_bore_62_ram_hold(sigFromSrams_bore_62_ram_hold),
        .sigFromSrams_bore_62_ram_bypass(sigFromSrams_bore_62_ram_bypass),
        .sigFromSrams_bore_62_ram_bp_clken(sigFromSrams_bore_62_ram_bp_clken),
        .sigFromSrams_bore_62_ram_aux_clk(sigFromSrams_bore_62_ram_aux_clk),
        .sigFromSrams_bore_62_ram_aux_ckbp(sigFromSrams_bore_62_ram_aux_ckbp),
        .sigFromSrams_bore_62_ram_mcp_hold(sigFromSrams_bore_62_ram_mcp_hold),
        .sigFromSrams_bore_62_cgen(sigFromSrams_bore_62_cgen),
        .sigFromSrams_bore_63_ram_hold(sigFromSrams_bore_63_ram_hold),
        .sigFromSrams_bore_63_ram_bypass(sigFromSrams_bore_63_ram_bypass),
        .sigFromSrams_bore_63_ram_bp_clken(sigFromSrams_bore_63_ram_bp_clken),
        .sigFromSrams_bore_63_ram_aux_clk(sigFromSrams_bore_63_ram_aux_clk),
        .sigFromSrams_bore_63_ram_aux_ckbp(sigFromSrams_bore_63_ram_aux_ckbp),
        .sigFromSrams_bore_63_ram_mcp_hold(sigFromSrams_bore_63_ram_mcp_hold),
        .sigFromSrams_bore_63_cgen(sigFromSrams_bore_63_cgen),
        .sigFromSrams_bore_64_ram_hold(sigFromSrams_bore_64_ram_hold),
        .sigFromSrams_bore_64_ram_bypass(sigFromSrams_bore_64_ram_bypass),
        .sigFromSrams_bore_64_ram_bp_clken(sigFromSrams_bore_64_ram_bp_clken),
        .sigFromSrams_bore_64_ram_aux_clk(sigFromSrams_bore_64_ram_aux_clk),
        .sigFromSrams_bore_64_ram_aux_ckbp(sigFromSrams_bore_64_ram_aux_ckbp),
        .sigFromSrams_bore_64_ram_mcp_hold(sigFromSrams_bore_64_ram_mcp_hold),
        .sigFromSrams_bore_64_cgen(sigFromSrams_bore_64_cgen),
        .sigFromSrams_bore_65_ram_hold(sigFromSrams_bore_65_ram_hold),
        .sigFromSrams_bore_65_ram_bypass(sigFromSrams_bore_65_ram_bypass),
        .sigFromSrams_bore_65_ram_bp_clken(sigFromSrams_bore_65_ram_bp_clken),
        .sigFromSrams_bore_65_ram_aux_clk(sigFromSrams_bore_65_ram_aux_clk),
        .sigFromSrams_bore_65_ram_aux_ckbp(sigFromSrams_bore_65_ram_aux_ckbp),
        .sigFromSrams_bore_65_ram_mcp_hold(sigFromSrams_bore_65_ram_mcp_hold),
        .sigFromSrams_bore_65_cgen(sigFromSrams_bore_65_cgen),
        .sigFromSrams_bore_66_ram_hold(sigFromSrams_bore_66_ram_hold),
        .sigFromSrams_bore_66_ram_bypass(sigFromSrams_bore_66_ram_bypass),
        .sigFromSrams_bore_66_ram_bp_clken(sigFromSrams_bore_66_ram_bp_clken),
        .sigFromSrams_bore_66_ram_aux_clk(sigFromSrams_bore_66_ram_aux_clk),
        .sigFromSrams_bore_66_ram_aux_ckbp(sigFromSrams_bore_66_ram_aux_ckbp),
        .sigFromSrams_bore_66_ram_mcp_hold(sigFromSrams_bore_66_ram_mcp_hold),
        .sigFromSrams_bore_66_cgen(sigFromSrams_bore_66_cgen),
        .sigFromSrams_bore_67_ram_hold(sigFromSrams_bore_67_ram_hold),
        .sigFromSrams_bore_67_ram_bypass(sigFromSrams_bore_67_ram_bypass),
        .sigFromSrams_bore_67_ram_bp_clken(sigFromSrams_bore_67_ram_bp_clken),
        .sigFromSrams_bore_67_ram_aux_clk(sigFromSrams_bore_67_ram_aux_clk),
        .sigFromSrams_bore_67_ram_aux_ckbp(sigFromSrams_bore_67_ram_aux_ckbp),
        .sigFromSrams_bore_67_ram_mcp_hold(sigFromSrams_bore_67_ram_mcp_hold),
        .sigFromSrams_bore_67_cgen(sigFromSrams_bore_67_cgen),
        .sigFromSrams_bore_68_ram_hold(sigFromSrams_bore_68_ram_hold),
        .sigFromSrams_bore_68_ram_bypass(sigFromSrams_bore_68_ram_bypass),
        .sigFromSrams_bore_68_ram_bp_clken(sigFromSrams_bore_68_ram_bp_clken),
        .sigFromSrams_bore_68_ram_aux_clk(sigFromSrams_bore_68_ram_aux_clk),
        .sigFromSrams_bore_68_ram_aux_ckbp(sigFromSrams_bore_68_ram_aux_ckbp),
        .sigFromSrams_bore_68_ram_mcp_hold(sigFromSrams_bore_68_ram_mcp_hold),
        .sigFromSrams_bore_68_cgen(sigFromSrams_bore_68_cgen),
        .sigFromSrams_bore_69_ram_hold(sigFromSrams_bore_69_ram_hold),
        .sigFromSrams_bore_69_ram_bypass(sigFromSrams_bore_69_ram_bypass),
        .sigFromSrams_bore_69_ram_bp_clken(sigFromSrams_bore_69_ram_bp_clken),
        .sigFromSrams_bore_69_ram_aux_clk(sigFromSrams_bore_69_ram_aux_clk),
        .sigFromSrams_bore_69_ram_aux_ckbp(sigFromSrams_bore_69_ram_aux_ckbp),
        .sigFromSrams_bore_69_ram_mcp_hold(sigFromSrams_bore_69_ram_mcp_hold),
        .sigFromSrams_bore_69_cgen(sigFromSrams_bore_69_cgen),
        .sigFromSrams_bore_70_ram_hold(sigFromSrams_bore_70_ram_hold),
        .sigFromSrams_bore_70_ram_bypass(sigFromSrams_bore_70_ram_bypass),
        .sigFromSrams_bore_70_ram_bp_clken(sigFromSrams_bore_70_ram_bp_clken),
        .sigFromSrams_bore_70_ram_aux_clk(sigFromSrams_bore_70_ram_aux_clk),
        .sigFromSrams_bore_70_ram_aux_ckbp(sigFromSrams_bore_70_ram_aux_ckbp),
        .sigFromSrams_bore_70_ram_mcp_hold(sigFromSrams_bore_70_ram_mcp_hold),
        .sigFromSrams_bore_70_cgen(sigFromSrams_bore_70_cgen),
        .sigFromSrams_bore_71_ram_hold(sigFromSrams_bore_71_ram_hold),
        .sigFromSrams_bore_71_ram_bypass(sigFromSrams_bore_71_ram_bypass),
        .sigFromSrams_bore_71_ram_bp_clken(sigFromSrams_bore_71_ram_bp_clken),
        .sigFromSrams_bore_71_ram_aux_clk(sigFromSrams_bore_71_ram_aux_clk),
        .sigFromSrams_bore_71_ram_aux_ckbp(sigFromSrams_bore_71_ram_aux_ckbp),
        .sigFromSrams_bore_71_ram_mcp_hold(sigFromSrams_bore_71_ram_mcp_hold),
        .sigFromSrams_bore_71_cgen(sigFromSrams_bore_71_cgen),
        .sigFromSrams_bore_72_ram_hold(sigFromSrams_bore_72_ram_hold),
        .sigFromSrams_bore_72_ram_bypass(sigFromSrams_bore_72_ram_bypass),
        .sigFromSrams_bore_72_ram_bp_clken(sigFromSrams_bore_72_ram_bp_clken),
        .sigFromSrams_bore_72_ram_aux_clk(sigFromSrams_bore_72_ram_aux_clk),
        .sigFromSrams_bore_72_ram_aux_ckbp(sigFromSrams_bore_72_ram_aux_ckbp),
        .sigFromSrams_bore_72_ram_mcp_hold(sigFromSrams_bore_72_ram_mcp_hold),
        .sigFromSrams_bore_72_cgen(sigFromSrams_bore_72_cgen),
        .sigFromSrams_bore_73_ram_hold(sigFromSrams_bore_73_ram_hold),
        .sigFromSrams_bore_73_ram_bypass(sigFromSrams_bore_73_ram_bypass),
        .sigFromSrams_bore_73_ram_bp_clken(sigFromSrams_bore_73_ram_bp_clken),
        .sigFromSrams_bore_73_ram_aux_clk(sigFromSrams_bore_73_ram_aux_clk),
        .sigFromSrams_bore_73_ram_aux_ckbp(sigFromSrams_bore_73_ram_aux_ckbp),
        .sigFromSrams_bore_73_ram_mcp_hold(sigFromSrams_bore_73_ram_mcp_hold),
        .sigFromSrams_bore_73_cgen(sigFromSrams_bore_73_cgen),
        .sigFromSrams_bore_74_ram_hold(sigFromSrams_bore_74_ram_hold),
        .sigFromSrams_bore_74_ram_bypass(sigFromSrams_bore_74_ram_bypass),
        .sigFromSrams_bore_74_ram_bp_clken(sigFromSrams_bore_74_ram_bp_clken),
        .sigFromSrams_bore_74_ram_aux_clk(sigFromSrams_bore_74_ram_aux_clk),
        .sigFromSrams_bore_74_ram_aux_ckbp(sigFromSrams_bore_74_ram_aux_ckbp),
        .sigFromSrams_bore_74_ram_mcp_hold(sigFromSrams_bore_74_ram_mcp_hold),
        .sigFromSrams_bore_74_cgen(sigFromSrams_bore_74_cgen),
        .sigFromSrams_bore_75_ram_hold(sigFromSrams_bore_75_ram_hold),
        .sigFromSrams_bore_75_ram_bypass(sigFromSrams_bore_75_ram_bypass),
        .sigFromSrams_bore_75_ram_bp_clken(sigFromSrams_bore_75_ram_bp_clken),
        .sigFromSrams_bore_75_ram_aux_clk(sigFromSrams_bore_75_ram_aux_clk),
        .sigFromSrams_bore_75_ram_aux_ckbp(sigFromSrams_bore_75_ram_aux_ckbp),
        .sigFromSrams_bore_75_ram_mcp_hold(sigFromSrams_bore_75_ram_mcp_hold),
        .sigFromSrams_bore_75_cgen(sigFromSrams_bore_75_cgen),
        .sigFromSrams_bore_76_ram_hold(sigFromSrams_bore_76_ram_hold),
        .sigFromSrams_bore_76_ram_bypass(sigFromSrams_bore_76_ram_bypass),
        .sigFromSrams_bore_76_ram_bp_clken(sigFromSrams_bore_76_ram_bp_clken),
        .sigFromSrams_bore_76_ram_aux_clk(sigFromSrams_bore_76_ram_aux_clk),
        .sigFromSrams_bore_76_ram_aux_ckbp(sigFromSrams_bore_76_ram_aux_ckbp),
        .sigFromSrams_bore_76_ram_mcp_hold(sigFromSrams_bore_76_ram_mcp_hold),
        .sigFromSrams_bore_76_cgen(sigFromSrams_bore_76_cgen),
        .sigFromSrams_bore_77_ram_hold(sigFromSrams_bore_77_ram_hold),
        .sigFromSrams_bore_77_ram_bypass(sigFromSrams_bore_77_ram_bypass),
        .sigFromSrams_bore_77_ram_bp_clken(sigFromSrams_bore_77_ram_bp_clken),
        .sigFromSrams_bore_77_ram_aux_clk(sigFromSrams_bore_77_ram_aux_clk),
        .sigFromSrams_bore_77_ram_aux_ckbp(sigFromSrams_bore_77_ram_aux_ckbp),
        .sigFromSrams_bore_77_ram_mcp_hold(sigFromSrams_bore_77_ram_mcp_hold),
        .sigFromSrams_bore_77_cgen(sigFromSrams_bore_77_cgen),
        .sigFromSrams_bore_78_ram_hold(sigFromSrams_bore_78_ram_hold),
        .sigFromSrams_bore_78_ram_bypass(sigFromSrams_bore_78_ram_bypass),
        .sigFromSrams_bore_78_ram_bp_clken(sigFromSrams_bore_78_ram_bp_clken),
        .sigFromSrams_bore_78_ram_aux_clk(sigFromSrams_bore_78_ram_aux_clk),
        .sigFromSrams_bore_78_ram_aux_ckbp(sigFromSrams_bore_78_ram_aux_ckbp),
        .sigFromSrams_bore_78_ram_mcp_hold(sigFromSrams_bore_78_ram_mcp_hold),
        .sigFromSrams_bore_78_cgen(sigFromSrams_bore_78_cgen),
        .sigFromSrams_bore_79_ram_hold(sigFromSrams_bore_79_ram_hold),
        .sigFromSrams_bore_79_ram_bypass(sigFromSrams_bore_79_ram_bypass),
        .sigFromSrams_bore_79_ram_bp_clken(sigFromSrams_bore_79_ram_bp_clken),
        .sigFromSrams_bore_79_ram_aux_clk(sigFromSrams_bore_79_ram_aux_clk),
        .sigFromSrams_bore_79_ram_aux_ckbp(sigFromSrams_bore_79_ram_aux_ckbp),
        .sigFromSrams_bore_79_ram_mcp_hold(sigFromSrams_bore_79_ram_mcp_hold),
        .sigFromSrams_bore_79_cgen(sigFromSrams_bore_79_cgen),
        .sigFromSrams_bore_80_ram_hold(sigFromSrams_bore_80_ram_hold),
        .sigFromSrams_bore_80_ram_bypass(sigFromSrams_bore_80_ram_bypass),
        .sigFromSrams_bore_80_ram_bp_clken(sigFromSrams_bore_80_ram_bp_clken),
        .sigFromSrams_bore_80_ram_aux_clk(sigFromSrams_bore_80_ram_aux_clk),
        .sigFromSrams_bore_80_ram_aux_ckbp(sigFromSrams_bore_80_ram_aux_ckbp),
        .sigFromSrams_bore_80_ram_mcp_hold(sigFromSrams_bore_80_ram_mcp_hold),
        .sigFromSrams_bore_80_cgen(sigFromSrams_bore_80_cgen),
        .sigFromSrams_bore_81_ram_hold(sigFromSrams_bore_81_ram_hold),
        .sigFromSrams_bore_81_ram_bypass(sigFromSrams_bore_81_ram_bypass),
        .sigFromSrams_bore_81_ram_bp_clken(sigFromSrams_bore_81_ram_bp_clken),
        .sigFromSrams_bore_81_ram_aux_clk(sigFromSrams_bore_81_ram_aux_clk),
        .sigFromSrams_bore_81_ram_aux_ckbp(sigFromSrams_bore_81_ram_aux_ckbp),
        .sigFromSrams_bore_81_ram_mcp_hold(sigFromSrams_bore_81_ram_mcp_hold),
        .sigFromSrams_bore_81_cgen(sigFromSrams_bore_81_cgen),
        .sigFromSrams_bore_82_ram_hold(sigFromSrams_bore_82_ram_hold),
        .sigFromSrams_bore_82_ram_bypass(sigFromSrams_bore_82_ram_bypass),
        .sigFromSrams_bore_82_ram_bp_clken(sigFromSrams_bore_82_ram_bp_clken),
        .sigFromSrams_bore_82_ram_aux_clk(sigFromSrams_bore_82_ram_aux_clk),
        .sigFromSrams_bore_82_ram_aux_ckbp(sigFromSrams_bore_82_ram_aux_ckbp),
        .sigFromSrams_bore_82_ram_mcp_hold(sigFromSrams_bore_82_ram_mcp_hold),
        .sigFromSrams_bore_82_cgen(sigFromSrams_bore_82_cgen),
        .sigFromSrams_bore_83_ram_hold(sigFromSrams_bore_83_ram_hold),
        .sigFromSrams_bore_83_ram_bypass(sigFromSrams_bore_83_ram_bypass),
        .sigFromSrams_bore_83_ram_bp_clken(sigFromSrams_bore_83_ram_bp_clken),
        .sigFromSrams_bore_83_ram_aux_clk(sigFromSrams_bore_83_ram_aux_clk),
        .sigFromSrams_bore_83_ram_aux_ckbp(sigFromSrams_bore_83_ram_aux_ckbp),
        .sigFromSrams_bore_83_ram_mcp_hold(sigFromSrams_bore_83_ram_mcp_hold),
        .sigFromSrams_bore_83_cgen(sigFromSrams_bore_83_cgen),
        .sigFromSrams_bore_84_ram_hold(sigFromSrams_bore_84_ram_hold),
        .sigFromSrams_bore_84_ram_bypass(sigFromSrams_bore_84_ram_bypass),
        .sigFromSrams_bore_84_ram_bp_clken(sigFromSrams_bore_84_ram_bp_clken),
        .sigFromSrams_bore_84_ram_aux_clk(sigFromSrams_bore_84_ram_aux_clk),
        .sigFromSrams_bore_84_ram_aux_ckbp(sigFromSrams_bore_84_ram_aux_ckbp),
        .sigFromSrams_bore_84_ram_mcp_hold(sigFromSrams_bore_84_ram_mcp_hold),
        .sigFromSrams_bore_84_cgen(sigFromSrams_bore_84_cgen),
        .sigFromSrams_bore_85_ram_hold(sigFromSrams_bore_85_ram_hold),
        .sigFromSrams_bore_85_ram_bypass(sigFromSrams_bore_85_ram_bypass),
        .sigFromSrams_bore_85_ram_bp_clken(sigFromSrams_bore_85_ram_bp_clken),
        .sigFromSrams_bore_85_ram_aux_clk(sigFromSrams_bore_85_ram_aux_clk),
        .sigFromSrams_bore_85_ram_aux_ckbp(sigFromSrams_bore_85_ram_aux_ckbp),
        .sigFromSrams_bore_85_ram_mcp_hold(sigFromSrams_bore_85_ram_mcp_hold),
        .sigFromSrams_bore_85_cgen(sigFromSrams_bore_85_cgen),
        .sigFromSrams_bore_86_ram_hold(sigFromSrams_bore_86_ram_hold),
        .sigFromSrams_bore_86_ram_bypass(sigFromSrams_bore_86_ram_bypass),
        .sigFromSrams_bore_86_ram_bp_clken(sigFromSrams_bore_86_ram_bp_clken),
        .sigFromSrams_bore_86_ram_aux_clk(sigFromSrams_bore_86_ram_aux_clk),
        .sigFromSrams_bore_86_ram_aux_ckbp(sigFromSrams_bore_86_ram_aux_ckbp),
        .sigFromSrams_bore_86_ram_mcp_hold(sigFromSrams_bore_86_ram_mcp_hold),
        .sigFromSrams_bore_86_cgen(sigFromSrams_bore_86_cgen),
        .sigFromSrams_bore_87_ram_hold(sigFromSrams_bore_87_ram_hold),
        .sigFromSrams_bore_87_ram_bypass(sigFromSrams_bore_87_ram_bypass),
        .sigFromSrams_bore_87_ram_bp_clken(sigFromSrams_bore_87_ram_bp_clken),
        .sigFromSrams_bore_87_ram_aux_clk(sigFromSrams_bore_87_ram_aux_clk),
        .sigFromSrams_bore_87_ram_aux_ckbp(sigFromSrams_bore_87_ram_aux_ckbp),
        .sigFromSrams_bore_87_ram_mcp_hold(sigFromSrams_bore_87_ram_mcp_hold),
        .sigFromSrams_bore_87_cgen(sigFromSrams_bore_87_cgen),
        .sigFromSrams_bore_88_ram_hold(sigFromSrams_bore_88_ram_hold),
        .sigFromSrams_bore_88_ram_bypass(sigFromSrams_bore_88_ram_bypass),
        .sigFromSrams_bore_88_ram_bp_clken(sigFromSrams_bore_88_ram_bp_clken),
        .sigFromSrams_bore_88_ram_aux_clk(sigFromSrams_bore_88_ram_aux_clk),
        .sigFromSrams_bore_88_ram_aux_ckbp(sigFromSrams_bore_88_ram_aux_ckbp),
        .sigFromSrams_bore_88_ram_mcp_hold(sigFromSrams_bore_88_ram_mcp_hold),
        .sigFromSrams_bore_88_cgen(sigFromSrams_bore_88_cgen),
        .sigFromSrams_bore_89_ram_hold(sigFromSrams_bore_89_ram_hold),
        .sigFromSrams_bore_89_ram_bypass(sigFromSrams_bore_89_ram_bypass),
        .sigFromSrams_bore_89_ram_bp_clken(sigFromSrams_bore_89_ram_bp_clken),
        .sigFromSrams_bore_89_ram_aux_clk(sigFromSrams_bore_89_ram_aux_clk),
        .sigFromSrams_bore_89_ram_aux_ckbp(sigFromSrams_bore_89_ram_aux_ckbp),
        .sigFromSrams_bore_89_ram_mcp_hold(sigFromSrams_bore_89_ram_mcp_hold),
        .sigFromSrams_bore_89_cgen(sigFromSrams_bore_89_cgen),
        .sigFromSrams_bore_90_ram_hold(sigFromSrams_bore_90_ram_hold),
        .sigFromSrams_bore_90_ram_bypass(sigFromSrams_bore_90_ram_bypass),
        .sigFromSrams_bore_90_ram_bp_clken(sigFromSrams_bore_90_ram_bp_clken),
        .sigFromSrams_bore_90_ram_aux_clk(sigFromSrams_bore_90_ram_aux_clk),
        .sigFromSrams_bore_90_ram_aux_ckbp(sigFromSrams_bore_90_ram_aux_ckbp),
        .sigFromSrams_bore_90_ram_mcp_hold(sigFromSrams_bore_90_ram_mcp_hold),
        .sigFromSrams_bore_90_cgen(sigFromSrams_bore_90_cgen),
        .sigFromSrams_bore_91_ram_hold(sigFromSrams_bore_91_ram_hold),
        .sigFromSrams_bore_91_ram_bypass(sigFromSrams_bore_91_ram_bypass),
        .sigFromSrams_bore_91_ram_bp_clken(sigFromSrams_bore_91_ram_bp_clken),
        .sigFromSrams_bore_91_ram_aux_clk(sigFromSrams_bore_91_ram_aux_clk),
        .sigFromSrams_bore_91_ram_aux_ckbp(sigFromSrams_bore_91_ram_aux_ckbp),
        .sigFromSrams_bore_91_ram_mcp_hold(sigFromSrams_bore_91_ram_mcp_hold),
        .sigFromSrams_bore_91_cgen(sigFromSrams_bore_91_cgen),
        .sigFromSrams_bore_92_ram_hold(sigFromSrams_bore_92_ram_hold),
        .sigFromSrams_bore_92_ram_bypass(sigFromSrams_bore_92_ram_bypass),
        .sigFromSrams_bore_92_ram_bp_clken(sigFromSrams_bore_92_ram_bp_clken),
        .sigFromSrams_bore_92_ram_aux_clk(sigFromSrams_bore_92_ram_aux_clk),
        .sigFromSrams_bore_92_ram_aux_ckbp(sigFromSrams_bore_92_ram_aux_ckbp),
        .sigFromSrams_bore_92_ram_mcp_hold(sigFromSrams_bore_92_ram_mcp_hold),
        .sigFromSrams_bore_92_cgen(sigFromSrams_bore_92_cgen),
        .sigFromSrams_bore_93_ram_hold(sigFromSrams_bore_93_ram_hold),
        .sigFromSrams_bore_93_ram_bypass(sigFromSrams_bore_93_ram_bypass),
        .sigFromSrams_bore_93_ram_bp_clken(sigFromSrams_bore_93_ram_bp_clken),
        .sigFromSrams_bore_93_ram_aux_clk(sigFromSrams_bore_93_ram_aux_clk),
        .sigFromSrams_bore_93_ram_aux_ckbp(sigFromSrams_bore_93_ram_aux_ckbp),
        .sigFromSrams_bore_93_ram_mcp_hold(sigFromSrams_bore_93_ram_mcp_hold),
        .sigFromSrams_bore_93_cgen(sigFromSrams_bore_93_cgen),
        .sigFromSrams_bore_94_ram_hold(sigFromSrams_bore_94_ram_hold),
        .sigFromSrams_bore_94_ram_bypass(sigFromSrams_bore_94_ram_bypass),
        .sigFromSrams_bore_94_ram_bp_clken(sigFromSrams_bore_94_ram_bp_clken),
        .sigFromSrams_bore_94_ram_aux_clk(sigFromSrams_bore_94_ram_aux_clk),
        .sigFromSrams_bore_94_ram_aux_ckbp(sigFromSrams_bore_94_ram_aux_ckbp),
        .sigFromSrams_bore_94_ram_mcp_hold(sigFromSrams_bore_94_ram_mcp_hold),
        .sigFromSrams_bore_94_cgen(sigFromSrams_bore_94_cgen),
        .sigFromSrams_bore_95_ram_hold(sigFromSrams_bore_95_ram_hold),
        .sigFromSrams_bore_95_ram_bypass(sigFromSrams_bore_95_ram_bypass),
        .sigFromSrams_bore_95_ram_bp_clken(sigFromSrams_bore_95_ram_bp_clken),
        .sigFromSrams_bore_95_ram_aux_clk(sigFromSrams_bore_95_ram_aux_clk),
        .sigFromSrams_bore_95_ram_aux_ckbp(sigFromSrams_bore_95_ram_aux_ckbp),
        .sigFromSrams_bore_95_ram_mcp_hold(sigFromSrams_bore_95_ram_mcp_hold),
        .sigFromSrams_bore_95_cgen(sigFromSrams_bore_95_cgen),
        .sigFromSrams_bore_96_ram_hold(sigFromSrams_bore_96_ram_hold),
        .sigFromSrams_bore_96_ram_bypass(sigFromSrams_bore_96_ram_bypass),
        .sigFromSrams_bore_96_ram_bp_clken(sigFromSrams_bore_96_ram_bp_clken),
        .sigFromSrams_bore_96_ram_aux_clk(sigFromSrams_bore_96_ram_aux_clk),
        .sigFromSrams_bore_96_ram_aux_ckbp(sigFromSrams_bore_96_ram_aux_ckbp),
        .sigFromSrams_bore_96_ram_mcp_hold(sigFromSrams_bore_96_ram_mcp_hold),
        .sigFromSrams_bore_96_cgen(sigFromSrams_bore_96_cgen),
        .sigFromSrams_bore_97_ram_hold(sigFromSrams_bore_97_ram_hold),
        .sigFromSrams_bore_97_ram_bypass(sigFromSrams_bore_97_ram_bypass),
        .sigFromSrams_bore_97_ram_bp_clken(sigFromSrams_bore_97_ram_bp_clken),
        .sigFromSrams_bore_97_ram_aux_clk(sigFromSrams_bore_97_ram_aux_clk),
        .sigFromSrams_bore_97_ram_aux_ckbp(sigFromSrams_bore_97_ram_aux_ckbp),
        .sigFromSrams_bore_97_ram_mcp_hold(sigFromSrams_bore_97_ram_mcp_hold),
        .sigFromSrams_bore_97_cgen(sigFromSrams_bore_97_cgen),
        .sigFromSrams_bore_98_ram_hold(sigFromSrams_bore_98_ram_hold),
        .sigFromSrams_bore_98_ram_bypass(sigFromSrams_bore_98_ram_bypass),
        .sigFromSrams_bore_98_ram_bp_clken(sigFromSrams_bore_98_ram_bp_clken),
        .sigFromSrams_bore_98_ram_aux_clk(sigFromSrams_bore_98_ram_aux_clk),
        .sigFromSrams_bore_98_ram_aux_ckbp(sigFromSrams_bore_98_ram_aux_ckbp),
        .sigFromSrams_bore_98_ram_mcp_hold(sigFromSrams_bore_98_ram_mcp_hold),
        .sigFromSrams_bore_98_cgen(sigFromSrams_bore_98_cgen),
        .sigFromSrams_bore_99_ram_hold(sigFromSrams_bore_99_ram_hold),
        .sigFromSrams_bore_99_ram_bypass(sigFromSrams_bore_99_ram_bypass),
        .sigFromSrams_bore_99_ram_bp_clken(sigFromSrams_bore_99_ram_bp_clken),
        .sigFromSrams_bore_99_ram_aux_clk(sigFromSrams_bore_99_ram_aux_clk),
        .sigFromSrams_bore_99_ram_aux_ckbp(sigFromSrams_bore_99_ram_aux_ckbp),
        .sigFromSrams_bore_99_ram_mcp_hold(sigFromSrams_bore_99_ram_mcp_hold),
        .sigFromSrams_bore_99_cgen(sigFromSrams_bore_99_cgen),
        .sigFromSrams_bore_100_ram_hold(sigFromSrams_bore_100_ram_hold),
        .sigFromSrams_bore_100_ram_bypass(sigFromSrams_bore_100_ram_bypass),
        .sigFromSrams_bore_100_ram_bp_clken(sigFromSrams_bore_100_ram_bp_clken),
        .sigFromSrams_bore_100_ram_aux_clk(sigFromSrams_bore_100_ram_aux_clk),
        .sigFromSrams_bore_100_ram_aux_ckbp(sigFromSrams_bore_100_ram_aux_ckbp),
        .sigFromSrams_bore_100_ram_mcp_hold(sigFromSrams_bore_100_ram_mcp_hold),
        .sigFromSrams_bore_100_cgen(sigFromSrams_bore_100_cgen),
        .sigFromSrams_bore_101_ram_hold(sigFromSrams_bore_101_ram_hold),
        .sigFromSrams_bore_101_ram_bypass(sigFromSrams_bore_101_ram_bypass),
        .sigFromSrams_bore_101_ram_bp_clken(sigFromSrams_bore_101_ram_bp_clken),
        .sigFromSrams_bore_101_ram_aux_clk(sigFromSrams_bore_101_ram_aux_clk),
        .sigFromSrams_bore_101_ram_aux_ckbp(sigFromSrams_bore_101_ram_aux_ckbp),
        .sigFromSrams_bore_101_ram_mcp_hold(sigFromSrams_bore_101_ram_mcp_hold),
        .sigFromSrams_bore_101_cgen(sigFromSrams_bore_101_cgen),
        .sigFromSrams_bore_102_ram_hold(sigFromSrams_bore_102_ram_hold),
        .sigFromSrams_bore_102_ram_bypass(sigFromSrams_bore_102_ram_bypass),
        .sigFromSrams_bore_102_ram_bp_clken(sigFromSrams_bore_102_ram_bp_clken),
        .sigFromSrams_bore_102_ram_aux_clk(sigFromSrams_bore_102_ram_aux_clk),
        .sigFromSrams_bore_102_ram_aux_ckbp(sigFromSrams_bore_102_ram_aux_ckbp),
        .sigFromSrams_bore_102_ram_mcp_hold(sigFromSrams_bore_102_ram_mcp_hold),
        .sigFromSrams_bore_102_cgen(sigFromSrams_bore_102_cgen),
        .sigFromSrams_bore_103_ram_hold(sigFromSrams_bore_103_ram_hold),
        .sigFromSrams_bore_103_ram_bypass(sigFromSrams_bore_103_ram_bypass),
        .sigFromSrams_bore_103_ram_bp_clken(sigFromSrams_bore_103_ram_bp_clken),
        .sigFromSrams_bore_103_ram_aux_clk(sigFromSrams_bore_103_ram_aux_clk),
        .sigFromSrams_bore_103_ram_aux_ckbp(sigFromSrams_bore_103_ram_aux_ckbp),
        .sigFromSrams_bore_103_ram_mcp_hold(sigFromSrams_bore_103_ram_mcp_hold),
        .sigFromSrams_bore_103_cgen(sigFromSrams_bore_103_cgen),
        .sigFromSrams_bore_104_ram_hold(sigFromSrams_bore_104_ram_hold),
        .sigFromSrams_bore_104_ram_bypass(sigFromSrams_bore_104_ram_bypass),
        .sigFromSrams_bore_104_ram_bp_clken(sigFromSrams_bore_104_ram_bp_clken),
        .sigFromSrams_bore_104_ram_aux_clk(sigFromSrams_bore_104_ram_aux_clk),
        .sigFromSrams_bore_104_ram_aux_ckbp(sigFromSrams_bore_104_ram_aux_ckbp),
        .sigFromSrams_bore_104_ram_mcp_hold(sigFromSrams_bore_104_ram_mcp_hold),
        .sigFromSrams_bore_104_cgen(sigFromSrams_bore_104_cgen),
        .sigFromSrams_bore_105_ram_hold(sigFromSrams_bore_105_ram_hold),
        .sigFromSrams_bore_105_ram_bypass(sigFromSrams_bore_105_ram_bypass),
        .sigFromSrams_bore_105_ram_bp_clken(sigFromSrams_bore_105_ram_bp_clken),
        .sigFromSrams_bore_105_ram_aux_clk(sigFromSrams_bore_105_ram_aux_clk),
        .sigFromSrams_bore_105_ram_aux_ckbp(sigFromSrams_bore_105_ram_aux_ckbp),
        .sigFromSrams_bore_105_ram_mcp_hold(sigFromSrams_bore_105_ram_mcp_hold),
        .sigFromSrams_bore_105_cgen(sigFromSrams_bore_105_cgen),
        .sigFromSrams_bore_106_ram_hold(sigFromSrams_bore_106_ram_hold),
        .sigFromSrams_bore_106_ram_bypass(sigFromSrams_bore_106_ram_bypass),
        .sigFromSrams_bore_106_ram_bp_clken(sigFromSrams_bore_106_ram_bp_clken),
        .sigFromSrams_bore_106_ram_aux_clk(sigFromSrams_bore_106_ram_aux_clk),
        .sigFromSrams_bore_106_ram_aux_ckbp(sigFromSrams_bore_106_ram_aux_ckbp),
        .sigFromSrams_bore_106_ram_mcp_hold(sigFromSrams_bore_106_ram_mcp_hold),
        .sigFromSrams_bore_106_cgen(sigFromSrams_bore_106_cgen),
        .sigFromSrams_bore_107_ram_hold(sigFromSrams_bore_107_ram_hold),
        .sigFromSrams_bore_107_ram_bypass(sigFromSrams_bore_107_ram_bypass),
        .sigFromSrams_bore_107_ram_bp_clken(sigFromSrams_bore_107_ram_bp_clken),
        .sigFromSrams_bore_107_ram_aux_clk(sigFromSrams_bore_107_ram_aux_clk),
        .sigFromSrams_bore_107_ram_aux_ckbp(sigFromSrams_bore_107_ram_aux_ckbp),
        .sigFromSrams_bore_107_ram_mcp_hold(sigFromSrams_bore_107_ram_mcp_hold),
        .sigFromSrams_bore_107_cgen(sigFromSrams_bore_107_cgen),
        .sigFromSrams_bore_108_ram_hold(sigFromSrams_bore_108_ram_hold),
        .sigFromSrams_bore_108_ram_bypass(sigFromSrams_bore_108_ram_bypass),
        .sigFromSrams_bore_108_ram_bp_clken(sigFromSrams_bore_108_ram_bp_clken),
        .sigFromSrams_bore_108_ram_aux_clk(sigFromSrams_bore_108_ram_aux_clk),
        .sigFromSrams_bore_108_ram_aux_ckbp(sigFromSrams_bore_108_ram_aux_ckbp),
        .sigFromSrams_bore_108_ram_mcp_hold(sigFromSrams_bore_108_ram_mcp_hold),
        .sigFromSrams_bore_108_cgen(sigFromSrams_bore_108_cgen),
        .sigFromSrams_bore_109_ram_hold(sigFromSrams_bore_109_ram_hold),
        .sigFromSrams_bore_109_ram_bypass(sigFromSrams_bore_109_ram_bypass),
        .sigFromSrams_bore_109_ram_bp_clken(sigFromSrams_bore_109_ram_bp_clken),
        .sigFromSrams_bore_109_ram_aux_clk(sigFromSrams_bore_109_ram_aux_clk),
        .sigFromSrams_bore_109_ram_aux_ckbp(sigFromSrams_bore_109_ram_aux_ckbp),
        .sigFromSrams_bore_109_ram_mcp_hold(sigFromSrams_bore_109_ram_mcp_hold),
        .sigFromSrams_bore_109_cgen(sigFromSrams_bore_109_cgen),
        .sigFromSrams_bore_110_ram_hold(sigFromSrams_bore_110_ram_hold),
        .sigFromSrams_bore_110_ram_bypass(sigFromSrams_bore_110_ram_bypass),
        .sigFromSrams_bore_110_ram_bp_clken(sigFromSrams_bore_110_ram_bp_clken),
        .sigFromSrams_bore_110_ram_aux_clk(sigFromSrams_bore_110_ram_aux_clk),
        .sigFromSrams_bore_110_ram_aux_ckbp(sigFromSrams_bore_110_ram_aux_ckbp),
        .sigFromSrams_bore_110_ram_mcp_hold(sigFromSrams_bore_110_ram_mcp_hold),
        .sigFromSrams_bore_110_cgen(sigFromSrams_bore_110_cgen),
        .sigFromSrams_bore_111_ram_hold(sigFromSrams_bore_111_ram_hold),
        .sigFromSrams_bore_111_ram_bypass(sigFromSrams_bore_111_ram_bypass),
        .sigFromSrams_bore_111_ram_bp_clken(sigFromSrams_bore_111_ram_bp_clken),
        .sigFromSrams_bore_111_ram_aux_clk(sigFromSrams_bore_111_ram_aux_clk),
        .sigFromSrams_bore_111_ram_aux_ckbp(sigFromSrams_bore_111_ram_aux_ckbp),
        .sigFromSrams_bore_111_ram_mcp_hold(sigFromSrams_bore_111_ram_mcp_hold),
        .sigFromSrams_bore_111_cgen(sigFromSrams_bore_111_cgen),
        .sigFromSrams_bore_112_ram_hold(sigFromSrams_bore_112_ram_hold),
        .sigFromSrams_bore_112_ram_bypass(sigFromSrams_bore_112_ram_bypass),
        .sigFromSrams_bore_112_ram_bp_clken(sigFromSrams_bore_112_ram_bp_clken),
        .sigFromSrams_bore_112_ram_aux_clk(sigFromSrams_bore_112_ram_aux_clk),
        .sigFromSrams_bore_112_ram_aux_ckbp(sigFromSrams_bore_112_ram_aux_ckbp),
        .sigFromSrams_bore_112_ram_mcp_hold(sigFromSrams_bore_112_ram_mcp_hold),
        .sigFromSrams_bore_112_cgen(sigFromSrams_bore_112_cgen),
        .sigFromSrams_bore_113_ram_hold(sigFromSrams_bore_113_ram_hold),
        .sigFromSrams_bore_113_ram_bypass(sigFromSrams_bore_113_ram_bypass),
        .sigFromSrams_bore_113_ram_bp_clken(sigFromSrams_bore_113_ram_bp_clken),
        .sigFromSrams_bore_113_ram_aux_clk(sigFromSrams_bore_113_ram_aux_clk),
        .sigFromSrams_bore_113_ram_aux_ckbp(sigFromSrams_bore_113_ram_aux_ckbp),
        .sigFromSrams_bore_113_ram_mcp_hold(sigFromSrams_bore_113_ram_mcp_hold),
        .sigFromSrams_bore_113_cgen(sigFromSrams_bore_113_cgen),
        .sigFromSrams_bore_114_ram_hold(sigFromSrams_bore_114_ram_hold),
        .sigFromSrams_bore_114_ram_bypass(sigFromSrams_bore_114_ram_bypass),
        .sigFromSrams_bore_114_ram_bp_clken(sigFromSrams_bore_114_ram_bp_clken),
        .sigFromSrams_bore_114_ram_aux_clk(sigFromSrams_bore_114_ram_aux_clk),
        .sigFromSrams_bore_114_ram_aux_ckbp(sigFromSrams_bore_114_ram_aux_ckbp),
        .sigFromSrams_bore_114_ram_mcp_hold(sigFromSrams_bore_114_ram_mcp_hold),
        .sigFromSrams_bore_114_cgen(sigFromSrams_bore_114_cgen),
        .sigFromSrams_bore_115_ram_hold(sigFromSrams_bore_115_ram_hold),
        .sigFromSrams_bore_115_ram_bypass(sigFromSrams_bore_115_ram_bypass),
        .sigFromSrams_bore_115_ram_bp_clken(sigFromSrams_bore_115_ram_bp_clken),
        .sigFromSrams_bore_115_ram_aux_clk(sigFromSrams_bore_115_ram_aux_clk),
        .sigFromSrams_bore_115_ram_aux_ckbp(sigFromSrams_bore_115_ram_aux_ckbp),
        .sigFromSrams_bore_115_ram_mcp_hold(sigFromSrams_bore_115_ram_mcp_hold),
        .sigFromSrams_bore_115_cgen(sigFromSrams_bore_115_cgen),
        .sigFromSrams_bore_116_ram_hold(sigFromSrams_bore_116_ram_hold),
        .sigFromSrams_bore_116_ram_bypass(sigFromSrams_bore_116_ram_bypass),
        .sigFromSrams_bore_116_ram_bp_clken(sigFromSrams_bore_116_ram_bp_clken),
        .sigFromSrams_bore_116_ram_aux_clk(sigFromSrams_bore_116_ram_aux_clk),
        .sigFromSrams_bore_116_ram_aux_ckbp(sigFromSrams_bore_116_ram_aux_ckbp),
        .sigFromSrams_bore_116_ram_mcp_hold(sigFromSrams_bore_116_ram_mcp_hold),
        .sigFromSrams_bore_116_cgen(sigFromSrams_bore_116_cgen),
        .sigFromSrams_bore_117_ram_hold(sigFromSrams_bore_117_ram_hold),
        .sigFromSrams_bore_117_ram_bypass(sigFromSrams_bore_117_ram_bypass),
        .sigFromSrams_bore_117_ram_bp_clken(sigFromSrams_bore_117_ram_bp_clken),
        .sigFromSrams_bore_117_ram_aux_clk(sigFromSrams_bore_117_ram_aux_clk),
        .sigFromSrams_bore_117_ram_aux_ckbp(sigFromSrams_bore_117_ram_aux_ckbp),
        .sigFromSrams_bore_117_ram_mcp_hold(sigFromSrams_bore_117_ram_mcp_hold),
        .sigFromSrams_bore_117_cgen(sigFromSrams_bore_117_cgen),
        .sigFromSrams_bore_118_ram_hold(sigFromSrams_bore_118_ram_hold),
        .sigFromSrams_bore_118_ram_bypass(sigFromSrams_bore_118_ram_bypass),
        .sigFromSrams_bore_118_ram_bp_clken(sigFromSrams_bore_118_ram_bp_clken),
        .sigFromSrams_bore_118_ram_aux_clk(sigFromSrams_bore_118_ram_aux_clk),
        .sigFromSrams_bore_118_ram_aux_ckbp(sigFromSrams_bore_118_ram_aux_ckbp),
        .sigFromSrams_bore_118_ram_mcp_hold(sigFromSrams_bore_118_ram_mcp_hold),
        .sigFromSrams_bore_118_cgen(sigFromSrams_bore_118_cgen),
        .sigFromSrams_bore_119_ram_hold(sigFromSrams_bore_119_ram_hold),
        .sigFromSrams_bore_119_ram_bypass(sigFromSrams_bore_119_ram_bypass),
        .sigFromSrams_bore_119_ram_bp_clken(sigFromSrams_bore_119_ram_bp_clken),
        .sigFromSrams_bore_119_ram_aux_clk(sigFromSrams_bore_119_ram_aux_clk),
        .sigFromSrams_bore_119_ram_aux_ckbp(sigFromSrams_bore_119_ram_aux_ckbp),
        .sigFromSrams_bore_119_ram_mcp_hold(sigFromSrams_bore_119_ram_mcp_hold),
        .sigFromSrams_bore_119_cgen(sigFromSrams_bore_119_cgen),
        .sigFromSrams_bore_120_ram_hold(sigFromSrams_bore_120_ram_hold),
        .sigFromSrams_bore_120_ram_bypass(sigFromSrams_bore_120_ram_bypass),
        .sigFromSrams_bore_120_ram_bp_clken(sigFromSrams_bore_120_ram_bp_clken),
        .sigFromSrams_bore_120_ram_aux_clk(sigFromSrams_bore_120_ram_aux_clk),
        .sigFromSrams_bore_120_ram_aux_ckbp(sigFromSrams_bore_120_ram_aux_ckbp),
        .sigFromSrams_bore_120_ram_mcp_hold(sigFromSrams_bore_120_ram_mcp_hold),
        .sigFromSrams_bore_120_cgen(sigFromSrams_bore_120_cgen),
        .sigFromSrams_bore_121_ram_hold(sigFromSrams_bore_121_ram_hold),
        .sigFromSrams_bore_121_ram_bypass(sigFromSrams_bore_121_ram_bypass),
        .sigFromSrams_bore_121_ram_bp_clken(sigFromSrams_bore_121_ram_bp_clken),
        .sigFromSrams_bore_121_ram_aux_clk(sigFromSrams_bore_121_ram_aux_clk),
        .sigFromSrams_bore_121_ram_aux_ckbp(sigFromSrams_bore_121_ram_aux_ckbp),
        .sigFromSrams_bore_121_ram_mcp_hold(sigFromSrams_bore_121_ram_mcp_hold),
        .sigFromSrams_bore_121_cgen(sigFromSrams_bore_121_cgen),
        .sigFromSrams_bore_122_ram_hold(sigFromSrams_bore_122_ram_hold),
        .sigFromSrams_bore_122_ram_bypass(sigFromSrams_bore_122_ram_bypass),
        .sigFromSrams_bore_122_ram_bp_clken(sigFromSrams_bore_122_ram_bp_clken),
        .sigFromSrams_bore_122_ram_aux_clk(sigFromSrams_bore_122_ram_aux_clk),
        .sigFromSrams_bore_122_ram_aux_ckbp(sigFromSrams_bore_122_ram_aux_ckbp),
        .sigFromSrams_bore_122_ram_mcp_hold(sigFromSrams_bore_122_ram_mcp_hold),
        .sigFromSrams_bore_122_cgen(sigFromSrams_bore_122_cgen),
        .sigFromSrams_bore_123_ram_hold(sigFromSrams_bore_123_ram_hold),
        .sigFromSrams_bore_123_ram_bypass(sigFromSrams_bore_123_ram_bypass),
        .sigFromSrams_bore_123_ram_bp_clken(sigFromSrams_bore_123_ram_bp_clken),
        .sigFromSrams_bore_123_ram_aux_clk(sigFromSrams_bore_123_ram_aux_clk),
        .sigFromSrams_bore_123_ram_aux_ckbp(sigFromSrams_bore_123_ram_aux_ckbp),
        .sigFromSrams_bore_123_ram_mcp_hold(sigFromSrams_bore_123_ram_mcp_hold),
        .sigFromSrams_bore_123_cgen(sigFromSrams_bore_123_cgen),
        .sigFromSrams_bore_124_ram_hold(sigFromSrams_bore_124_ram_hold),
        .sigFromSrams_bore_124_ram_bypass(sigFromSrams_bore_124_ram_bypass),
        .sigFromSrams_bore_124_ram_bp_clken(sigFromSrams_bore_124_ram_bp_clken),
        .sigFromSrams_bore_124_ram_aux_clk(sigFromSrams_bore_124_ram_aux_clk),
        .sigFromSrams_bore_124_ram_aux_ckbp(sigFromSrams_bore_124_ram_aux_ckbp),
        .sigFromSrams_bore_124_ram_mcp_hold(sigFromSrams_bore_124_ram_mcp_hold),
        .sigFromSrams_bore_124_cgen(sigFromSrams_bore_124_cgen),
        .sigFromSrams_bore_125_ram_hold(sigFromSrams_bore_125_ram_hold),
        .sigFromSrams_bore_125_ram_bypass(sigFromSrams_bore_125_ram_bypass),
        .sigFromSrams_bore_125_ram_bp_clken(sigFromSrams_bore_125_ram_bp_clken),
        .sigFromSrams_bore_125_ram_aux_clk(sigFromSrams_bore_125_ram_aux_clk),
        .sigFromSrams_bore_125_ram_aux_ckbp(sigFromSrams_bore_125_ram_aux_ckbp),
        .sigFromSrams_bore_125_ram_mcp_hold(sigFromSrams_bore_125_ram_mcp_hold),
        .sigFromSrams_bore_125_cgen(sigFromSrams_bore_125_cgen),
        .sigFromSrams_bore_126_ram_hold(sigFromSrams_bore_126_ram_hold),
        .sigFromSrams_bore_126_ram_bypass(sigFromSrams_bore_126_ram_bypass),
        .sigFromSrams_bore_126_ram_bp_clken(sigFromSrams_bore_126_ram_bp_clken),
        .sigFromSrams_bore_126_ram_aux_clk(sigFromSrams_bore_126_ram_aux_clk),
        .sigFromSrams_bore_126_ram_aux_ckbp(sigFromSrams_bore_126_ram_aux_ckbp),
        .sigFromSrams_bore_126_ram_mcp_hold(sigFromSrams_bore_126_ram_mcp_hold),
        .sigFromSrams_bore_126_cgen(sigFromSrams_bore_126_cgen),
        .sigFromSrams_bore_127_ram_hold(sigFromSrams_bore_127_ram_hold),
        .sigFromSrams_bore_127_ram_bypass(sigFromSrams_bore_127_ram_bypass),
        .sigFromSrams_bore_127_ram_bp_clken(sigFromSrams_bore_127_ram_bp_clken),
        .sigFromSrams_bore_127_ram_aux_clk(sigFromSrams_bore_127_ram_aux_clk),
        .sigFromSrams_bore_127_ram_aux_ckbp(sigFromSrams_bore_127_ram_aux_ckbp),
        .sigFromSrams_bore_127_ram_mcp_hold(sigFromSrams_bore_127_ram_mcp_hold),
        .sigFromSrams_bore_127_cgen(sigFromSrams_bore_127_cgen),
        .sigFromSrams_bore_128_ram_hold(sigFromSrams_bore_128_ram_hold),
        .sigFromSrams_bore_128_ram_bypass(sigFromSrams_bore_128_ram_bypass),
        .sigFromSrams_bore_128_ram_bp_clken(sigFromSrams_bore_128_ram_bp_clken),
        .sigFromSrams_bore_128_ram_aux_clk(sigFromSrams_bore_128_ram_aux_clk),
        .sigFromSrams_bore_128_ram_aux_ckbp(sigFromSrams_bore_128_ram_aux_ckbp),
        .sigFromSrams_bore_128_ram_mcp_hold(sigFromSrams_bore_128_ram_mcp_hold),
        .sigFromSrams_bore_128_cgen(sigFromSrams_bore_128_cgen),
        .sigFromSrams_bore_129_ram_hold(sigFromSrams_bore_129_ram_hold),
        .sigFromSrams_bore_129_ram_bypass(sigFromSrams_bore_129_ram_bypass),
        .sigFromSrams_bore_129_ram_bp_clken(sigFromSrams_bore_129_ram_bp_clken),
        .sigFromSrams_bore_129_ram_aux_clk(sigFromSrams_bore_129_ram_aux_clk),
        .sigFromSrams_bore_129_ram_aux_ckbp(sigFromSrams_bore_129_ram_aux_ckbp),
        .sigFromSrams_bore_129_ram_mcp_hold(sigFromSrams_bore_129_ram_mcp_hold),
        .sigFromSrams_bore_129_cgen(sigFromSrams_bore_129_cgen),
        .sigFromSrams_bore_130_ram_hold(sigFromSrams_bore_130_ram_hold),
        .sigFromSrams_bore_130_ram_bypass(sigFromSrams_bore_130_ram_bypass),
        .sigFromSrams_bore_130_ram_bp_clken(sigFromSrams_bore_130_ram_bp_clken),
        .sigFromSrams_bore_130_ram_aux_clk(sigFromSrams_bore_130_ram_aux_clk),
        .sigFromSrams_bore_130_ram_aux_ckbp(sigFromSrams_bore_130_ram_aux_ckbp),
        .sigFromSrams_bore_130_ram_mcp_hold(sigFromSrams_bore_130_ram_mcp_hold),
        .sigFromSrams_bore_130_cgen(sigFromSrams_bore_130_cgen),
        .sigFromSrams_bore_131_ram_hold(sigFromSrams_bore_131_ram_hold),
        .sigFromSrams_bore_131_ram_bypass(sigFromSrams_bore_131_ram_bypass),
        .sigFromSrams_bore_131_ram_bp_clken(sigFromSrams_bore_131_ram_bp_clken),
        .sigFromSrams_bore_131_ram_aux_clk(sigFromSrams_bore_131_ram_aux_clk),
        .sigFromSrams_bore_131_ram_aux_ckbp(sigFromSrams_bore_131_ram_aux_ckbp),
        .sigFromSrams_bore_131_ram_mcp_hold(sigFromSrams_bore_131_ram_mcp_hold),
        .sigFromSrams_bore_131_cgen(sigFromSrams_bore_131_cgen),
        .sigFromSrams_bore_132_ram_hold(sigFromSrams_bore_132_ram_hold),
        .sigFromSrams_bore_132_ram_bypass(sigFromSrams_bore_132_ram_bypass),
        .sigFromSrams_bore_132_ram_bp_clken(sigFromSrams_bore_132_ram_bp_clken),
        .sigFromSrams_bore_132_ram_aux_clk(sigFromSrams_bore_132_ram_aux_clk),
        .sigFromSrams_bore_132_ram_aux_ckbp(sigFromSrams_bore_132_ram_aux_ckbp),
        .sigFromSrams_bore_132_ram_mcp_hold(sigFromSrams_bore_132_ram_mcp_hold),
        .sigFromSrams_bore_132_cgen(sigFromSrams_bore_132_cgen),
        .sigFromSrams_bore_133_ram_hold(sigFromSrams_bore_133_ram_hold),
        .sigFromSrams_bore_133_ram_bypass(sigFromSrams_bore_133_ram_bypass),
        .sigFromSrams_bore_133_ram_bp_clken(sigFromSrams_bore_133_ram_bp_clken),
        .sigFromSrams_bore_133_ram_aux_clk(sigFromSrams_bore_133_ram_aux_clk),
        .sigFromSrams_bore_133_ram_aux_ckbp(sigFromSrams_bore_133_ram_aux_ckbp),
        .sigFromSrams_bore_133_ram_mcp_hold(sigFromSrams_bore_133_ram_mcp_hold),
        .sigFromSrams_bore_133_cgen(sigFromSrams_bore_133_cgen),
        .sigFromSrams_bore_134_ram_hold(sigFromSrams_bore_134_ram_hold),
        .sigFromSrams_bore_134_ram_bypass(sigFromSrams_bore_134_ram_bypass),
        .sigFromSrams_bore_134_ram_bp_clken(sigFromSrams_bore_134_ram_bp_clken),
        .sigFromSrams_bore_134_ram_aux_clk(sigFromSrams_bore_134_ram_aux_clk),
        .sigFromSrams_bore_134_ram_aux_ckbp(sigFromSrams_bore_134_ram_aux_ckbp),
        .sigFromSrams_bore_134_ram_mcp_hold(sigFromSrams_bore_134_ram_mcp_hold),
        .sigFromSrams_bore_134_cgen(sigFromSrams_bore_134_cgen),
        .sigFromSrams_bore_135_ram_hold(sigFromSrams_bore_135_ram_hold),
        .sigFromSrams_bore_135_ram_bypass(sigFromSrams_bore_135_ram_bypass),
        .sigFromSrams_bore_135_ram_bp_clken(sigFromSrams_bore_135_ram_bp_clken),
        .sigFromSrams_bore_135_ram_aux_clk(sigFromSrams_bore_135_ram_aux_clk),
        .sigFromSrams_bore_135_ram_aux_ckbp(sigFromSrams_bore_135_ram_aux_ckbp),
        .sigFromSrams_bore_135_ram_mcp_hold(sigFromSrams_bore_135_ram_mcp_hold),
        .sigFromSrams_bore_135_cgen(sigFromSrams_bore_135_cgen),
        .sigFromSrams_bore_136_ram_hold(sigFromSrams_bore_136_ram_hold),
        .sigFromSrams_bore_136_ram_bypass(sigFromSrams_bore_136_ram_bypass),
        .sigFromSrams_bore_136_ram_bp_clken(sigFromSrams_bore_136_ram_bp_clken),
        .sigFromSrams_bore_136_ram_aux_clk(sigFromSrams_bore_136_ram_aux_clk),
        .sigFromSrams_bore_136_ram_aux_ckbp(sigFromSrams_bore_136_ram_aux_ckbp),
        .sigFromSrams_bore_136_ram_mcp_hold(sigFromSrams_bore_136_ram_mcp_hold),
        .sigFromSrams_bore_136_cgen(sigFromSrams_bore_136_cgen),
        .sigFromSrams_bore_137_ram_hold(sigFromSrams_bore_137_ram_hold),
        .sigFromSrams_bore_137_ram_bypass(sigFromSrams_bore_137_ram_bypass),
        .sigFromSrams_bore_137_ram_bp_clken(sigFromSrams_bore_137_ram_bp_clken),
        .sigFromSrams_bore_137_ram_aux_clk(sigFromSrams_bore_137_ram_aux_clk),
        .sigFromSrams_bore_137_ram_aux_ckbp(sigFromSrams_bore_137_ram_aux_ckbp),
        .sigFromSrams_bore_137_ram_mcp_hold(sigFromSrams_bore_137_ram_mcp_hold),
        .sigFromSrams_bore_137_cgen(sigFromSrams_bore_137_cgen),
        .sigFromSrams_bore_138_ram_hold(sigFromSrams_bore_138_ram_hold),
        .sigFromSrams_bore_138_ram_bypass(sigFromSrams_bore_138_ram_bypass),
        .sigFromSrams_bore_138_ram_bp_clken(sigFromSrams_bore_138_ram_bp_clken),
        .sigFromSrams_bore_138_ram_aux_clk(sigFromSrams_bore_138_ram_aux_clk),
        .sigFromSrams_bore_138_ram_aux_ckbp(sigFromSrams_bore_138_ram_aux_ckbp),
        .sigFromSrams_bore_138_ram_mcp_hold(sigFromSrams_bore_138_ram_mcp_hold),
        .sigFromSrams_bore_138_cgen(sigFromSrams_bore_138_cgen),
        .sigFromSrams_bore_139_ram_hold(sigFromSrams_bore_139_ram_hold),
        .sigFromSrams_bore_139_ram_bypass(sigFromSrams_bore_139_ram_bypass),
        .sigFromSrams_bore_139_ram_bp_clken(sigFromSrams_bore_139_ram_bp_clken),
        .sigFromSrams_bore_139_ram_aux_clk(sigFromSrams_bore_139_ram_aux_clk),
        .sigFromSrams_bore_139_ram_aux_ckbp(sigFromSrams_bore_139_ram_aux_ckbp),
        .sigFromSrams_bore_139_ram_mcp_hold(sigFromSrams_bore_139_ram_mcp_hold),
        .sigFromSrams_bore_139_cgen(sigFromSrams_bore_139_cgen),
        .sigFromSrams_bore_140_ram_hold(sigFromSrams_bore_140_ram_hold),
        .sigFromSrams_bore_140_ram_bypass(sigFromSrams_bore_140_ram_bypass),
        .sigFromSrams_bore_140_ram_bp_clken(sigFromSrams_bore_140_ram_bp_clken),
        .sigFromSrams_bore_140_ram_aux_clk(sigFromSrams_bore_140_ram_aux_clk),
        .sigFromSrams_bore_140_ram_aux_ckbp(sigFromSrams_bore_140_ram_aux_ckbp),
        .sigFromSrams_bore_140_ram_mcp_hold(sigFromSrams_bore_140_ram_mcp_hold),
        .sigFromSrams_bore_140_cgen(sigFromSrams_bore_140_cgen),
        .sigFromSrams_bore_141_ram_hold(sigFromSrams_bore_141_ram_hold),
        .sigFromSrams_bore_141_ram_bypass(sigFromSrams_bore_141_ram_bypass),
        .sigFromSrams_bore_141_ram_bp_clken(sigFromSrams_bore_141_ram_bp_clken),
        .sigFromSrams_bore_141_ram_aux_clk(sigFromSrams_bore_141_ram_aux_clk),
        .sigFromSrams_bore_141_ram_aux_ckbp(sigFromSrams_bore_141_ram_aux_ckbp),
        .sigFromSrams_bore_141_ram_mcp_hold(sigFromSrams_bore_141_ram_mcp_hold),
        .sigFromSrams_bore_141_cgen(sigFromSrams_bore_141_cgen),
        .sigFromSrams_bore_142_ram_hold(sigFromSrams_bore_142_ram_hold),
        .sigFromSrams_bore_142_ram_bypass(sigFromSrams_bore_142_ram_bypass),
        .sigFromSrams_bore_142_ram_bp_clken(sigFromSrams_bore_142_ram_bp_clken),
        .sigFromSrams_bore_142_ram_aux_clk(sigFromSrams_bore_142_ram_aux_clk),
        .sigFromSrams_bore_142_ram_aux_ckbp(sigFromSrams_bore_142_ram_aux_ckbp),
        .sigFromSrams_bore_142_ram_mcp_hold(sigFromSrams_bore_142_ram_mcp_hold),
        .sigFromSrams_bore_142_cgen(sigFromSrams_bore_142_cgen),
        .sigFromSrams_bore_143_ram_hold(sigFromSrams_bore_143_ram_hold),
        .sigFromSrams_bore_143_ram_bypass(sigFromSrams_bore_143_ram_bypass),
        .sigFromSrams_bore_143_ram_bp_clken(sigFromSrams_bore_143_ram_bp_clken),
        .sigFromSrams_bore_143_ram_aux_clk(sigFromSrams_bore_143_ram_aux_clk),
        .sigFromSrams_bore_143_ram_aux_ckbp(sigFromSrams_bore_143_ram_aux_ckbp),
        .sigFromSrams_bore_143_ram_mcp_hold(sigFromSrams_bore_143_ram_mcp_hold),
        .sigFromSrams_bore_143_cgen(sigFromSrams_bore_143_cgen)
    );

    assign io_toFtq_prediction_ready_o = io_toFtq_prediction_ready;
    assign s1_fire_o = dut.s1_fire;
    assign abtb_io_stageCtrl_s0_fire_probe_o = dut.abtb_io_stageCtrl_s0_fire_probe;

endmodule
